`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WPmBfcbnLEGINaiXUhLCWnGXhdziZJghPIpPpLU5FVDV1mIDHxz7UFnIbyhYnmPhoyoyKeThehqT
d6SZfjNs8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZQLIDsdxwDhnfh+8QKgBlqDUthjjX8VveYVLgIDucw1DWVXWofXQUABFgrMilan1yjE7aBoMSe++
01T9htQn3l9hMHNydDZ9QQ/cFtIuuvQJXs9Js84T4DilJn63BpHYGB5RmP4MJCacrL2JSNDzY+hG
RUFcwRxbj5FK0ImiTzY=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sCbOd2jalgBpJfH79h2qOT9EYfq69l68sKgObc8tSxcu89r1zJAfeqRUc60AKlstZq9MRiPG8moD
Z+wQbu97tOmHGUs5Q+P9jRTzR1YGxu4EWrL92ZTXJySrKtZjTgz68Gge2cRTtOtM4arEZgUAQrav
FRdisR/v/ro/KrXCS4U=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t2kui/PxWcDWEz2RkaNFrSqBGCaSFkcxUt9ZR1VEwKWu4YWAw0pDP4CHlmi6RL3wrPgqNm+JlVUf
fvYl2JMB2ZAiE0v0+Uhhta+IfKIO/OrK0tZGhfyK3lAr7x8QkG1pA7NfJ/8l+G8dw7ZaFCvCR34n
c5QhMSPcBEveqN4sBp/M7n9rmERmc7GtjX+vaPSRAGq3rLJFmCZs8GP9nu6UziJ4B1ThtIPgDrUl
uqZGrLY/uk5XMaezcsC/mQGMoAXL3IzE0uEeuUxCjaj4NMmaIGKXzqumOB+dOMV5Bhh7aCWH+ZSn
eqK5OFV0ItoUmvIpsNcgyGoQ9gqK0GS8SFNxOw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pAHup8Xf9xS9KRzEAWHDixdkKzJBOP87856UpROjyagDyFPHSWDGB5wCdx+cp2PKxh6EwzjfiQYw
bEP5Klayrlx8/NefyVw1WtNwCYzqFN/2NuHG/j3gKFSk3XMtsWUU9+YpVLkDpDF59dXTtp5Q5lvh
CEF/3TlGVgeGrS1agG5s7AgZBei7EQ9mHt74LzSMyrv1Hnk0pk7MnysYQDCglYgRXPoN4Q2euKgt
ZvtK1a57SKlRIUSc7mtkXanRLFX0WNH2YtLlSUo3CV719wgcUB4+yl9RJo+6u6G1TTcGoOHErngu
zduxtbFrxusro//gJEmgYq7hY3yCQTRROLIuMg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eHF0KjeEIXjNhmvZMvAKPRZTais/TzZ3YZ2ZVrLDBy2HUgd4Ux9YJlTeoPuUzJxh9IUobK+X5cLD
f5ufPEoR5uiNGe/+/Dw9q+jcKd5DH23jMK6vO9z+rAXbXqjTYIy67pDG06bIdh5yKi2IGpCrZfa+
kE6sfg1ZJYm6NDZ/GvXGdJ+oqewlcZ2jxdkj3E4+uotsGMrifG3ECwtHnIy2I+rvYj1smg7G7QTC
p3a8WF7aTqE2dWmIg9tJiCvwzON+f3W+q6Byy6AbIKWkBJhmtIls1iTwq1L1SdV2DhTJyINjbkfN
ifDV4PF6JK1wOdEdGRU2C4PqNYBwoF5wKf2NEA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 565792)
`protect data_block
4BZ1amLQ/23W4cc9WfV/IPSDcKabkp7d150n1e5ksDMSChMEEM5SIBUXGgCXqu+nOl2ihrk/wyq9
kBsWJPjI4bg2DI8/8mI977R34T+F+V6dcK5lT6wR1koC08dTtgPqThhYbs1ZqTWXlgTNYLUbd64f
+nz761jBJ5t6WK51xHhK4KONokoRrSmGA8A0EnIHCOvvXA7vUw0QSK6Bdy0ukNX/8K5XOeXn6sux
p+kqvl33U3SU+cakAlpzC1J6bmio9FdAo52pcCKkrjiwuv114V9d5MV9YcrDGIiAtMorRwZOIXNu
b+0vwEPrxp42kUpLyVAFY+al9ZoXu+HD0ubdJepnRECWFlTUTZ4uLW54fLJNn4lw7KQyiv/W/etC
RN9dyV66Dvf4CumOi0PfIWtq2gSMXx1R3ZeWmdcUM4wif+D4BgaE9iD92pf5tNTmXy9KfsxMN1/3
NiK7XPsvHxhsgHj4i54FfLqLXA/9rgNVEL9B62sQ72VnlZ5HoCPvZDwOC6aiXe55s6GdmLRmXFvb
09kwB5FzqDVgTX0IKQfFb670TVDtz/8MNI9PpZG3EhBljoW8D/8MxwfmWU19iw3aG6Iuaa5lGvWX
HZ0MkZWcN48ay3XeZYIx7M+FQ5SuZ/dgAD0tasL3vjy/2bQvJYJWK6fIP4avF6c6x2gAQz7oGbUB
cAP62TMsS+5Pa06VltWXmn/G8RlPEAYRsl3n9Gu32dUYo45v3hQVrD7lOHdxjz4cahN+XVlo8q6r
V34YDuFmMbhvK8WQ6Kg3UAwuOrNkP5Z2Ew6q7TZ0sT9wogbtLUZR//OGuMxrMvclKIJC4MuuAKbx
/MdnAr+8gfNNrACkWy/7eracu42sxFlElnNw0qb94DQrebJTgfJIQ3VmVtGkSA86zDFSgBC8/mI9
X4K5FPTOt62vLKanXUBj70/hLHBaqlt/ofgBS2Cb7OvOs5pxCTIQBD0JkzlQ45OMNIXxi7JnW9GG
CkIjYXHu4Y2VOs2HWqPDi/ZFiyHPm/4UkvtFI/VhJ8GB3XeL/tZqmCYDNx51Ovi/vmaM/sKQhJ4p
Haa7z2NukiyxHvCOyEo27ZRRQgmKNAXY/AbtWW78rRigORQpGbJupEbReCR26SsOzHTTciKjDbOJ
LVnasSjPqFZyhYyeVRVxDbLLOiVp9h9YjvIXJgqryCamU4y1GbafvSpkpCRmxGlr3T3rGRqsXhIS
dBDPw9p3yiLTcp1rCOr2s9mV0KjOMS6nKGzLbXaiRysdSPIJ0O8oQGY3RLGboQV6GQgtb9WLGyME
DmNiHUQEv6+AadSNjbjALFNLRnvXeh61D/dzWWM/eJWBqzTlfphk3zbHb0IW2gmN5UJxOhDNPrrE
P4SeUvsfKgI/DZiuovGI3gp/foDPpEo9/oCfb3jWYcQBd2TAnq27QSuDK7wyQeH5SxR3j1+LzkWu
SUB4dTT5sRjmObrHTl5Kd4Ut0v5hLVY3udoL6As6nNZcrMGmMA4UkBqLR0jBIKcCt5asJgT/Rw1b
MZ0ZqgK/beTMP9N8J+IF7CywBKfXSa34vffWwVqsfy9GvABO6w5YAtLpHBd8azwp4kYStyedxfxz
y1hx1ntIwX4Bw1LRGvPe70vWi6PwreS4vqq3Q2nacyF/neTyC6zxMbsOaJNCryYSikpfRac/zYRe
60mb3uA/9eqfmmzSitXwUHw+P8XRJ01qcQV9vAmO4I/BM0nb0l8o4rS9H1stX6O26uNK7T/9CXtW
uJ70w95s7H4MvH+1BTQoxq2KBta4XdxlriMmz7Q55ITCowcuG32tZnHYfTx45l/zpup69Laf7wUv
rWFGPlvn2tLOaFpY7qRY14RbuoP2h1cfR7jESzDHmIijQbJnxGe++RefGQ7E7ftc6RPYorC/ELoj
hgTgoB43muxVcT/UKMwKdRPO2KNLzLPyNEFLtIe7bWJZEZXOHF9JchOJ5OjE/pc0YRAHfGfYMhTf
eqwyj5j4ahq6LnK+8GGF9+pqc3UzkrhqY1PPeScQMJLyEJ/wPC9ELsIPm0s7PierSl56zqG48h3U
dEZL1j9MjVggUboudrLTDkIWHhjOrq2fyW3GCp02iCwlZR9eIUAyIos0wK6iMS7nXhQUv+rKaaWz
by/Xj0/OFqknGGqA0xiqyEZmtE4Xd3G0e7wGWKrXJxkqYFPaxCWsMAtdFTnFrE/w+onSqACWShce
3pGRoN6qsoCfjrzGrMgxrcsrRri6FqKmt1zY3LE3xY1g6R4B3ZisKpzG8m8aDSw9VZ/eeoCyuHYL
hfGvUeUneySZ8hM2U2/Qi3bJUCdVxgaGjrcZkXJeZ12Dxru8ha7ZVO7uzGjuK610kwBVOMTf2wwX
fIyncnbo+E2M2LvrXXUCtDhXn68U2bSFftmjwCYnE0kD2xn40CQn7jfQXqwE4oXPImi6q4CUgVYN
zM0bi7jiGcPtwJgG1R5gSlOMflfCApTdc42VbeCH2+6DH78cBYZ4uk3wWV89O8peE9hl0/9nN29z
cui+MH3xZ6mrh/OI2YJFJ+TNTZqjpOC6sU46dmSo4rUGfBC1FuIOzt0llsYOZff7uMNsDNtU7+/P
e2VOQoOwQ5OV9DBx1bQZXn5XZIC8qBDZFZexmMjAsNmLZEhxgAsOYZYgBUae7Nhjkk8vhx+DBap0
YLQtNDjpXWcxd0GEFp6cvNMx8MLQYeDD2tXZmoGeDPTIc5ST0ZCeC+aIdhXE+CxeeyfeWNSJLuts
WTIFuv8fXEz8JGWTMZ0fyL0e8r8YuGR6De4uq8IkWA6534R78yiO0ezJZL24WSgMow2jgHtsujll
ID4j98Jn1yId87YXd1ewElfBqeat9EeL5erVice9BeX9zexZYB3TC20Ci2ZYA+dK7Uv3dIjaFz6k
duchkczn8SOqFGiwlQkvbh/W68UKAPVMr4a4POPkVWOM+LNrixMvWCLXlttpih99mV8myN6mZBJd
oq7DJZ5ABvcPGN7KqXebTQHLaeDSiXhevYqIQVNTInblh8dte53rM+HrZeI9cjQtLTY5SQ0ROH39
2Al/uFg9/NvJdFJgLQGbbBpHP0o377BlOZhocmZJ0qOcELuGcFv22slNUNGH2aH8q3zvRdFEm2KY
3Jxn8EXtwVRz9rKKIMuEkonCtzGyFb2e3dhiZloTB1M9zlH2H9v0MCuqfFB+4XjOXldvQqdTAvA5
c4wk5CwmVrvXqVopwNbUNj3pCxvgzs2n8vy4Et6SiM0ztYgHCUZemS1sBq7K4SrrziZWvSN/zh/+
onehzT9Q0PYGYX9OPPwYzQ7VxqVWoaVbBKRIXLB52XO0s+gTLr97wIbssg1k9w3WHVbmnkWEW1lm
6VLOYJpbMfM4bf0erfaSmWZrkN4f4yEmrIM6xNZ6CMcIQPL+Y1Odl/4bEmcW+7BV+Ow8paOyPzQT
Fah5YEvwsPFSp/FTCBS4mcSQWLNhdj/tkcsvcT37Qm8DoFuQ/VkPjjacGxqZzRsyu0Xs+dCTnBxQ
Ae90/PRXF32j9xEHX7F0I0SLOY6s3xxFGXEnbH6GcAXfIyGRomxnLqsQ8n2x1HE6hq3V86ahIE9y
6kGnMdfh6re407W/aZs3vVkql/sAyVPdmi43srz1UiwlwwJ/rEJghceU0E5Yu99FaYbaVIhdbpEu
SwCajNv9c0hfWnJdRXeldzSorx9Rk5w3QzxZUArGdZWRWv5aXgQDKGzHWUZfhk/yVXAcZw0tJrfX
PieNZF8pLk+LgbSaf3ZVS8Ct6CqG5g62UOgpZDxsaUQ9q7OQ257IxRcs7bwd5UmDBl1WHu2ifjqP
toB5G1Wx6whOeGUCngs6Tsk3fu333ovW1HLfUEsgsb+jABmwLO/GokammDCNTU766iUZ9o7O6n9n
dlidjtKyHjSRwpZN4+xBrfcikl7F+Vx4yz1AyivAqlk2IO+2t78lo2o59wjRGY4ZAOYfS9wnTqG4
Mj4oUTZ30M3QRZnvdGqWfS23P3iHKa9hoDhknY0FrKhdTvlbmlEx7gNTzKuDZWDu+TAdbW5qF9/P
1ppUGuHoWN30SZ7ZnBl+ZhZr+Hu4TUoP8CY+u01mF1AHhefeUrnWdV8sBpz0y7Vzi3f7oSGRT1dM
+7HMX2K7kbimKT1SDPYzUHOJTvzPP4lEiH6GrWcQNkNxn1Shd0gITI8+iXUvY3V839C9z+M+CAzv
Y6S0xVIuZIgn2S0dt2md4xSeIGGrhPmrmk11DExPTOL2TPYCDwauv39JRxgzJi26cHzNf+VZDcw3
Z8SVR/6hf8sxv3cA1B1Cbav4R9Pi/6/hUBh9fXzxpZm0gcuGL5Ewvhd9uHBJUDozsL5DOQ/4HUJU
PkN1Mnqb+CSBPWXxLJl1g/PjCKMcbn/ucyCEiw5oUt1FWmcybu3GoAfy+ZRo8+2qWi9I+mWn++/v
0Oa1xV15chCT2yx0nrwrJHnotZPwyfheCYHIHqTtX+qHb79sn0uah37IxfmP+nfwex85Yq/u2tGK
yRT3s3VJKOcujm5Vhd8OmuRbI6pwmOa8i6b3VUYqh5YCYavx9P3YKDvBHogTaz2wSe9oJRm3/ZIA
YWpLH88iRU87w/43jdhT6rTOgfCEpc9WWxDYnYkzrzMsTKMO2HnCIsnqN/agz/j1Fyap1j/6vv6r
AYiDuB2+nsZmuauF7u/vEbUBpuKo63knQkQltFsoveMrenJBUUMipTbGfIYmnwMCHHELzMNm8eMv
zmwXDXQrD6lGlc1Pu4cKAO6oASpe/ifxLRviaipT8vKtW+hcxP0CqWeLriQ49eWMTfXx1zHRm3Jw
KWPqHHk8u+M+BvjDP0MkiKxU/RrvIJ0Pt7h9l2+KkOtishYtlhmx5EY4yH8G/SY2sIKA2XsduF/D
0BTe+CqCKMJxBy6wIljVGqEbpWnMi//s405frqxhDRgzV1p9jxffWLj3P/YidJ7KJkjV1/8i3MPB
hlzS88l4xnVlQ4frruZmKUJRXFbyIo9cgAg3p8gKNvSRelTnrtsDXftw8w0CrwGnpKpZ1a0f5nne
kNtGM5COIwFRu+v12IMusoD/mS/2eyhTb53H16sXbReFhnZthpySZ/kR/MhMdyMY1rYqIoYnKxMm
GYYwDbHoBrEsXEHpH6zCkW4+i8yjVa+KVRAiLOGi5NFgRZC1LkkjcurJ2sWHphFfGA41VoaehsuD
u6LTy5pAWlclmpoHIwo/ypFKrreRLkSa45C2Xjx9vgnkK988IB1dETXbKDk9634UOz4OBziialiq
hS8eD/uYaxhviyzo14hj73EERAinJ3Gh2K+exsj+bckDT28kgy9wxlJ5uc5R8V11LR/7qx5MuzXN
MD8ztRaS9fAMXn4CokX/1w02YrYr2bZrBBWryv3PKCdPG7s3PkBr7gTIlBwbtZv8wWgB4WsI+cY1
HH5Bv1pAEDho2KqkXeqSCvmxdqfU09oOFtt1JFBH3IhTk3ZXB86hAuQKApFqezhpOEG9LAalrUzT
9Qg+9G+q8TaOVWCQrACKumGxGKWd4GUIUFGZYHHupx/VCjiEfpq48WQwUtsCRbNfl1026DUQqtT3
/xoOA4sPQSRweMRZsxGHepXAF0eS3KJrzwB+dwS7MHpwteItygG/TgU5ecXTA8dacCDEcKajRfP+
7h9EDDj2gcmOVmISVE8PkEhyxU3KFmM+whzIxgvXpcB/afNfIEj9StPNHHTfbG/iXLEMIldQliDd
6MTow5T9XAkCQmFIQTwvI1ZYx9BMlk5YGeMlQIFJAMwt33raCSUmhWNGGMPGMJNtNDz/bkTk9XXw
TH97QzAYPiZ5VKo4NN6A0bHjlr32YAMcOJutbjF9X0T4Sy79ZjPzoXD1ZjXrL0XYKURLja1v+8N5
gL3HNZWrLaWsoVuSNV0dKCdOm9G+n4nfulXpMhvxXw28+39vcUFzh3gO/3ghI0NCXlgIiQtn/nu0
kVuyBJ+Veg60ugYaLAcfUUk67ZXaN64q6d1PNBGDaeTvF2rYWwZW5WCvik1FscEF6jBGh55vah6N
BQZf2wV2O8ftGB+2J6hAdwedgPLBzXo2WQEkRTC8qCW2GXq0DQohFqGkCEmK/elU/XOVSRx1Z1XH
gFEFT5dJ5lAmcXbRUv8IAsRB6FcmoYR3zeg+fkwWY1QUj+oAnMWkoUd1pW1mGKFtpYiyR1yc1FPH
c7KxoJZMWWUMfpdtBbc8mu7q+nuikc9TsF/3HABTiE+7RiL1tErU7iCJWMsezuCdXl3yKzwLfJib
5xjwhfBXInWBMelnSoKOCj4gWJMmt8Uxz2p3qVqBkhZ/54fuCYSHO6LV9l8lo6r5bHV9IUUaX1fH
52iM39SPBc316RFhmk+NydL4ja1Znw9Cvt5fVJT6Z493aoEwR90dpP0HE3xFKtx/L7w2OMt7gXBe
9pTHCnUfODul3P5RpUkYPd0Yqs9XGLdRb6jFOd3ZqXXjDDffY8YlTTGlJzWUeOv3iarGo1EUg3rc
VzBVSKrxZHbsxS+wTe/kAnlaSwkftu4BZ/qRpdKh3xJHW3g3YINOFIR68R+x1LE0YLABDQypTHPC
vVpZh9fVYrnRwKCF0QGqDCZweyuGDYhL2X0vGK6+r3/OoIseeL6S8pA6DzKbqN/62zL7HMroQ2Zk
yWQTzjHtozQr0Zd4Pp8Ev7FwTeH9kLcLZjhWnxS5AOuFjN2alUOCvHmhMhCWgOW45+tTYcoeefNQ
0Q+cv6Iqk2DX53XzLuKfbOjiffDxfYU0HUbwUwX7dZ+O/BGoUxBrHLQy8eAPl4GKuj3QXRIiiOPQ
UTyP6A02YhBwjDnMhw+qc0Fhe3xrclqL5pdk4LqSA4GR0Xezm2Z0n6uvIffKtMQvVmskLDyOB+Op
4vIvFtDmkV+G2ddx+4l1+7imUqdb88bdDjogO0xvOdwbZuAlVk2JSD0UWJtt+sRYzcpqN79qi0aM
98YRVNA9F774ed54cvYdgRI4NfdS+247IwJ73EKejlxCd6nPnP60kW4Pc0o3D1IQD7f8dWs+70Kz
qantK3hG+ce5Jbk599vKj/WKgv95JMu//ej7gNXsBQRhy0ukVe5hO9aSKB9N5NKFtgBzd/PQT0PP
OhkvsIs94FbCbcZLAtrcwfoTNzYN1knAKQUWxJWaTByTQ5iTAXtF0S2vIzSiA6XyBeyyH6l/ljpE
1veNAggOy0b+JtErRNnf8K42b8YLIFZ0whvTZ/qCn3NKMbxuviQFKc0/qQut4DzpIlIWZScQAJ5G
Kcbd/65izHf/HjgpwFLnLkaiToIttOto+GInXI5Qa7ABGrMqdmm5QJgev1Zsmg4OA27g/he+g9wG
ihO9Ha3Ju9f+QGJL3vpLD+VM4PMdLQSGwtrLkCc3t6fWunDAiRlOaCrgfi5IZJ1QGOH0W00lniJa
gCA5EZ1fuJNk22ZHEiMzo1ZIEaE77QjSxboanz00urOXX1Gb7ucn9VflQgUPrB1IugVvJnry29sr
gy1flnp6Czn3aE8QhQPgZXX+XS766FZffpeSobg7NKmUanwa38Sd0VbERtEHQq9RoJI/O7cpjcZE
2AUpeYROkodUsGfZxj74iCQzyIgXpy3TeQ4+iPNpa3/ohCVoR5Gk4QfqCPekcfbPBiCkIILhQlol
ODheDrfLzbr+yjeYzJqAwVPMy258aX1jI3XKGN3LmR+Qe5ervdWqeEN1S+lB4xJ38OWRAs8N1H3+
OcORKhDA6If+6a2QjC0ifrmbnoXLzDRYN7oybMx05tln3ySHBwCqi6TVFBXC/1L355Catq7iF6TL
7s69mL/rXCudn0Aq3VqlXOzPhdAMxM/Xf5wDTNo1Dy6onpLNtKlsu0W9qRo/5Dl9STPCRHemX7aB
AyprHEgrVW91f0eJA32Zkd0f87VqV09nSqurYv4kWDV+/853xdWprhersi6CL2YCt+L2cTIhMqmD
hiP1eKF2DBhGXSaU9TZ38hFAfc2yRgncL1r9JE879UKvexWNhSU1gt85bkJkD8GZpjmU8SJUMk+P
ec+kgBS+q8hs0UZmBZ5uYio7JSk2LRArpIb6RdP5mFCJimeH5WDpWNvY/hxyECV8plolC4Fp+BFi
ng/chqerDVyVdcI2qctoyjhVbmX0MPXesCCYKMa1awshVVMzbI+lkAzKeCkBvn+UhjB+N8v+3Fys
3Cao38H3uP2tI5PGDtTjT2n7SBAU8wK50qhjWK3agXdw0wxzsSFvqF76Ohzl/7XrBa154mNn7JG8
oMKMa56zoKhDxrFBR342154pRyPURyrFK60XjUpUoNaGQ5HUYH8CJcNm7Vm94jJdDdlBWU3zg0Jh
Z1mzdYxOyunbhqSoHvahBWCuCojJr4tCWwQTKHbS0BG5gf+4Cmd2B376Jd7ZzXckw6KkbrtotRui
OWfI3IKg3mNSGxqmt24+Fi8ZF/5dZrf/UKoq+IZ9uiZeZ82YbM2yNppA0v3+ZpbxnfRXE/eLryJT
8/UnOoEczaJSrpIwH/36S4Py6bfbGts4p6qKUjm/3a9iSFQotPGL7UlgZOba/keht6y7mfgvWu74
XKHCWpwQqrx1/2dY9RQrrwXmoF6xNYhHgYLCZPSShI1Q0i93JeDuM8+iv4MU/NKCEAvCNKvRLYyZ
hnizfmRmrEYJy7fOm2jpiIqHRls4ZTi60HruwbjSIMOMiEcUV+VDBx2OCwkL39+WoWCpNfKCrzCQ
4IP7a+DL1Xab4oB79mykgECYy2Cmm5u/xBFxuPg9JYKnpCnt4maEfWWfWrwmyF+3mLJPHCfkDlDU
rKn/eIWNgGc8xQGlOuAhDETjIjmLRPdi7Fi8Av5li66k1Sf8VYCaXjvGaXKk5Qqohy9Vtsx49ZZu
AyYthavA2NFp9YqIK4l0G74+cBPYQ4TRvcA5qdsaoXZjEnRQa48E3vqe8kMaVCHAkL11tRRiX2yl
RiExRoQwI/RtA9WU6YBrf66tJ+sxP8M8ofpOAGBljDmOUhLWS6OpHhir980ewgcf0ZRE/e8sHw3l
KBfplSk7za+eCyP+EyxOReOCQxeAyFGLIL9bMntj5nNK8z87gWn6A66aCW/zCcshaPSZCEZA34MT
BAsA4NdDsYGNKycH5n8lRAyPt9Y/xUQlEEJbtVMV5JzxF98MVKDO6CoJUCrUv8QorEobhTmRB2U5
XoyNb0zArl5RGdF2+MX+iOLtZV1tK9ERQM4SzDHu9brLbLCHm9prGXvId0OgjX5yfrgXDfN8k3Cz
ZzI8vfacxXRPZaAWY7jPDIWiTNC445kL2u7n0WDKPEuWzLSuDntVsR8bsteTJxT8gYytJ2liAj+w
4/k3xDY3grj1+5CxEzCZFv4qh+UItOfatuIGm4RBTEj6/f5rMAOwzfejTxygntbx5PD1faT5gwO/
WyBazg1xXujGq+lnm42DPxtEhT62aUkVinC/YzMl8oKbapibRNax7i2k4LrKvBKpkffFh2iCbJDx
7EzwewhUHlMEop0Qq489023Ola6DpwXvqbEHyFpslP3v0oXMBrT9Nhv5Y1xWJymBPC31TsxOqnGT
IH7/X7IQaKoaPB5LwFbS7P22ozL6TIVdZJpkJAfbBj5PfjNfA31WjYLpTU937P98KnG4fX1aR3QZ
Ku9E7Cd8ugK67UcXhVUWmZL7kuv1w9mLIxkLlMUXxitBDsNCPWbtaUQ8wckj1uCqmSl4iWjNYmn8
pJIJsiQxaiMWCXfFczy/xQaltSsq3ztE3mKt7gtbB4OpgJV2V8ur2eHRXdi4Q2a/IdRlfYKtkEa5
7e8nExqZJwo4tKjzntoLADmPLKD/p3oLIGuC3r5/jlkNTr93JSK5HP9HqhltEDcaHA3njS7NHbPX
uw6AwvNY5rDGGZJFtHiGZkmE6IYWypUVrTkecGPr41x+uSJ1r1BXMFfSs/pD0w2hKo3ExptlXDKF
nR0vjTOtIoBiERCToOPjy9gRdgD/wv6ol2/iEJsvI6fdG7jMv3aX/Dbcs7y9cLPgK2g65zJ0Xadv
XfE+cWPi8mK2L5s417e6K3O+dV3bWo714CigO4oG8gaFELPErw48I6Cr2XchRy91d2wjwH7kjeYM
1z+4QjAPSjhXUYvncxGLDLWUDhWwwoIrZTNz7n+AYxt3xSmYcsueU8p6oXWqERdlgbmldGDgMu3X
RLFms3rwUDeiTnr0EWAJ3e7GbfL4bP3yLgjCtwWHsIdO7NjV0WQ7mvgseDXt1eLaBT2Pj1arrUTK
EE23aAoMeSGfMECwZZjhcOuVogNlZ6LtejjP96xnBqsqGnnJqESJ3z8TiN9FkyQ8vfvkjypy9/Ho
hKUo+63wi3yau8vrjMbUbKcSZCG6/tyOrpj54QrBxOn/geoNyFozt31nEBVUKPuYlMV1P9D51+M+
aL7cqbky2wztPzJ1e3Uf5UXUNhG0/A9DWRclqCRqj4EfJVxBO2rh+nvFZLXBJskWOgqZJ9as4RdL
IwQgi8ndbQp2HuT6H71NcanSt8TP2ZTvpNE1LlVd8WHesWNa4/vG6uORv5c7KFn2TYEoOwL6K7Z2
cvb/9XzMdFcXMmZMr0TItpFlMVs+4AV9V8+dBlUK0J7KGaxPf61FiiZIapB6kvasLMzUwBD7Lqfy
lKmT6mnK9oZ8pOsQkaTEUqORNmEL+9yiCuUVnUTF1JKz7I1sDa1zKizbCvf47IsFnBfx0m7pjDQx
JU5PXruP2P6NShfCaxPg6L78th+dKsLEd2U9UUxFMK4UVsURxjH5i3E9VQp7u1g7wYn9X+H45JGU
M95iOD11Q9ksmgVdsYx46imCFVY2DIgnWTSyIjLCcTKzxuqEFz3tUrjcjgORl9XgEfwpSZqyidB4
O8dfxreit6jTQ3RpsCPVmxOoG4Dwkf15O92bVLhDCCJ34ZKtfur9HAJuMXieXzfpec7fSMz3viM8
BD1jB0kTbZbtK1obvJAg8caFKn2VkWmQeUG7wztkKt57YRy/jeykh0JE5ECdQXmec0TJLJ7dWEXz
Ic+AHQUG0fZUHQfT9bwNdqmx4R9fytKymF3D3JYBbQemNuJ3lrUDSwdFv4WFtuWVcMUbLge753LL
cKC7kASOnQJNtQlTxflsN6q4uoE0433R4C2hEzt+Sq3eN2qhHWKX6zSI8xJ+wnHgMGDWIMluVS3u
LdY7scNEMyWxv1ngfhwv1Egs0tZt53y2DRllJ5j1x6dI6hYshW8xVj2+g99V3HbFi7hgwN7iTQ8e
YcCJAysiP1RIB/Mic8S3UHF5G1+zXsLup8e4Lralf90/Z4TBCYa0ZBHQFfOZNDPoqgpOtR6V3afD
292yfOyD5QVXMRIFjBvsdOwLsPzvF+e3vR0j1hl7KkAC+/r5byClsBi9xbogV8Wbp6e9HRZVQfN5
RW/UCj92sTaP9dooeEZwSXh2YdX8p3fNWllCCfnCeqzdUTtmBcUouIKIfERARVXavO0mTPqdfRYw
xJXnoyuOYQz0U7wgTLN55SY/WXBaw/Bpw43BsOm8PReA2AnaIwo9lSR3YkrfDPty8CD6BXth9f20
lRKBaC8lFj3RFkZ0s/wBGl5LNRk4AeolRieqBdEMXNnJ7SY2BUgvxPFNPqDzbmHrQe1UxDH2gYtJ
33PviPHKeKDsKbMOFkPLAfRQga7xG9C615EkxP46HK2CMND+KT9kF8ZzWPzHuhEjCCLMSv/aZm3+
dTQBihlCSLewc80J+y5U3eYEu39BKcoobKPf0OLPqD/mCIGzSJwXknOdUAdbjeeKAt4EwBG46z9U
TslFC/4KTLt8s4lM41VjMOtGJGatdvdQv5oo5L+bbKEPTyo2J+JIJxkbDlyNicKml/IyJxDEB1om
isl3ZBNrqjnWwAg1dCxQFjAue//9cIpl4/srDEp/X1YfnY+4CXRKugbRYUBzU0WDv+x0sdy5ea/l
ZWm6Gp6shuK90DUimnrBddL+tTOnOObQFzrklQG/BkDKAYr8SmzOhY4xYH9SNcg3TMCtaq8tMFfo
wW4xPc2KNXMy0wWk0KUAOsNNQK2mTMnPmgrVTK2oiCPfHH2G1x5XV0DQNwcAU6o0+Jj9dAU72kJ1
r8juJjDaqE9QhN4OKe5DSDDyX9WQiS85DFF+DK4suhNCocsyojkNoyNPMCjUIiOwXOd0hm7KF+iR
qU1Ds/EUdFppooKFcO7D2IHux0gViyP/xupRHGa1VFrQ1TfkFFWYUDJUSNslhIowKlh+saMqc6vr
fKspsv+k7e8IahmOfcxevPR5T7IkEZYfcorNqLZ/zZYOZtnoNU9RPwCIU7wh9HdQ9jmXc9MPBBcV
oT965cuoefg1y5FL0TYYrOJDWwOjqZiXNQt8gca3TKAYM1QoIHUmcCowyMocS8++Szh5LpoJbzQJ
0RboziNNw4T/3LgHSg4B8MaFtfjzDKzgeA6Wb3t0n7vVo46hUrBj66odK0uOLy0kbobu8XOR83ic
cbe4Gh0JFx4qzLy1xVVs3oodAFTYQdaOy475dJKQ8ueNz4Otuhyn61nAjbSQD090Jh5LzutsFs3Y
B+LfpbOUVn17KZzA/XIXKF1fiPUYM7GuyFp0jbi+g8NCWKUULl3uJ2o+3zO8K/66GdDlFCUNs63e
3WpxBxwKqp1MwWPcl+JexOJOfFjLAeAC+T5sYU7DooINnr0vbjRhkJwON6IEe8DAfxh25Fdfm4m6
taWWv/6YjupaFqoQ6lgrrbu1QJCbrEfa/zEpzSff1gsVrdgf3Kg52OKxsos1yHCzonf7QWPm34aE
LJvxrnF9nu0ROuaoQhguPRnDfPiRX3csbhLyM6YPJSRVmHLd00oKh7pT5IExm23M/hKMX9ykI1T6
JP9Jlj8ibl/LFTXsPcwyLlniiU06ii7mMKhuSJI1wgbRb99UN9wK6+J9YAZ0XArKaFuOSC9SEK0i
BIlTq/Jyu+ZPv9mrl8jVsYeo/y7ini97Feup5LF4zhQbIeEysk7mYI6M/m2GXK2aqUR1z8DBp5un
gerfby/06TpGgf3BeWIh4GpnsCgBjv5m+5ygOQihoR/HrQAkt5ViQYEWnTAsK2Rf0o3p++2ak7kA
o1PiyGiQqysLGAX8a1zdNXI97aU3zTWQe6qYjTWk4yMBYm2frvPLV7RbmVGZvupa0mVC2R0wo2k8
9U4LEmIFm8DZ0VGwMLGdyy7ZeslOZ5difcbf35Xw/JotNeknM8qzKeAVvB7c8Jknioy3g7waEs9A
2S4Q4z9wvh+GTOD8SzjzGV1XbOsSqO1CBuejjU5LhBFRltcGng8sq7VM0B+FDlL0ax7Y+6XLAp/b
atPkVi11AqmqrPsPRofIcS5UytNIqbeylARX14P4fIUdc+XE1MZKGyYNkT+ObAmtXNlotL935ZE2
p8krqIyh6Va3gGTCdUbavorSMF3IEwjmZfXzGGq18eafGRA65OC6Y+EvdedUwY8lQrb4MNo7g8E/
zzrxferNJukWosUIkCzYKl2vXCA8svmN8xatRlhwSx34YLLluLBrUJSjrJGzOZwr6pP2xhODuvWy
NR2OdcDZVBIeimP0b3OF9eIVgcSFJXYMztmfjO7HZXdHNejwvVl4P3eEg/33wSyNonGhIFxbfJIj
9k1d5TjFo+bH9jw6ABxKxh8o460HypEYjjR7II76WiuVAf6kNTqTxQT1eu8EnY5ckxHkFSSMtemL
26thLb9NCvG7q6Ubi++Mt6LLAma57+1txiVySQq7ueDA5oPOb1aZE0MzWOvCf+Dl5bI1r8iKAmdn
0n2J9IN3LN3t887Y9b7uxl5uKy+Ec+pFBLU48yFT+CeRE5z9aD+I0zuAm6eYcvBD3dwTn9pCt0Ci
RVsKjM5SvTe9bVKjxO+Mt7Z74W2ZFZ1Gi0HWzLdCCe0BMB4KkiCzjasEoay3TRzf4Ld++j85SUvZ
2GWGdrQBdYpSCAzc3dOh7XNbv7znWY7CklYGj/8eKJ8ZMQk0H+FwnU7ogG0/E05pznWfIjnmVp20
BOTosPlPZjvd4d9ubi7C7MSGh5yKkOjnErH5NfptC8yoUO7UI2LszlMMSpQHARoHfsjUGq4OHCdE
+LevpikDOG2aDyjgOqVbZ1OJXNAUzloq2TKBPyhDCJLy+v87LJ7b5vgK1IW1DattAyQcdjl6doTl
WlGtSOHwrhGwQbWW/IOCWjxMq8R9FStdPpOyM8EKwZmRfMRKB2ivhuMA7XgkLPFCw/pW4gRKUjpd
fgG5RQnNts2aPu6Lmvv++fJnuZXIW+qpR7Yy1ojApYEq2mvXDdm3fkqI8YZowvFrLQkdE4nJbWW/
ESZEvFzT2xuguD9vqA+6woBcrSnzmV4/fneMs5T0apg/VFoIkyl207i3UM1xL7k2Z4JdG1K+faPK
R+qUvRtkBI3QNnrOjp23RCS5bhHBh2eDt3ykGacNZxE0CVz018ejAVyEiAId1TS81G8KzFV3h6B8
R1V2nEXwjQs9yqCkV4HrVO3g3cjbz0fcLKdgnhZgtJqRZBf51LbTRKbz/QIjVYQneZjq159vMZyL
kzoWt1EmoBoG79Nn9OB4TnNqcqVXP5q3UlwYbX/GbPHvHBEAqPwWblNJF2EGJiIPsBV00+eShxnh
IulqHukzXJUXmuY4IEyQzfFn+gybXQwJ04LR2GDAuN58Oxcci4WkNbZIQJmRCg97mq1wHETnk8av
HN7+shgPuSKcqYpdyc+o1ioHvcF1n9KttpNL4PdTxGoIvMl1p19RKQy/hvGQho0upHbguc/SShEq
Q1HNO5xQV6vJzRjVblUc7BiDEQopHDZj1WU/xnwYSz5sRXu6pgWY2+qa6lDit1zRqgOryyJEBCF8
ikCQ/vpzW2OjBQ7+wrzDdUPGqj9LIlG0vZsnzSislwrIl/jBxqtOqtLThMG044vjTaBSaIwrE1E/
mU7xJvu+IVHGid8p8WD3yEbdVL2BZMEZfkFDizNkOj5drkoyRRaimIM80iXxIW/5Y7otsYuA8AvZ
zCTfpVS+Gdnm+MoYw9xbcLL/M/AFs183Ip+bfC3ouWQuVakEhF9U4mHAXOvk93HcZoEie1T8l/BG
+uHOob/N1rqH4TaNUWhY1o74Wa4Yux/J9arc/il95TJhtLYaQMIbkSPOlpPJSeTyqCqfN9YKuupO
lGzuVX4N6f9UQs9jkbSl5qJ8LIJpKukpoOrS3gRpqnAVIFrSoPnoWt1czlC+tmyKZR2RCIiX7cik
jPC3ZQe1SitWTe0uaVwXUtYl0plStJ6Ks5/YPFBD5oSuBTpocW4/9P8QUtvitmlGLHWF0qVYN4Zw
Q9BMIhkbOZp61QbDLtzaxYQcKRv+mC85jntOxcaTUrBG+ic61rY+6JTF9Xo6kXhsF8iZcX+ZITh7
G9qJTqpokYRufd8gHGBFcvHwp5hC/hQg4i7kTKYZYR6ljf8PWGLfFB1nrSS8zC3sHjUAF+/juiWP
aUMjOxgHA+XsXCktq7H5yUOmkTh/e75USrL2tBKfPyw6jycVBClrICkeghe9l7KiOe4pAhCOJE7r
/5UHBUnNca130YifW0miF0/R9ecvFMc/wOgUA7/9PG13B4mpqxS7eJuT1rnophkUHYvHkhsgMf/V
3FYSAzQbSURdJOR0Yo5zcbL10j93ZIHoWzCbzLO28lJugal1Sh8ON8sXLnSQiR0jYqvSqSEtaVi0
1J7xaiMuqSez+4MTVf+I/NzdzS2q9flNU7Hb3xzZhyLz8ojHySZ/0TqnDhkrp8jdcPltANFCbBtg
FZ5A7o0p+qnnX3Nx+PAIBt3vh5Mozrz2dt9uyOEUgixj6M99Niu7TFD610a5R4K+37M13HGhGHnl
2c1pvDdloehJZRtWDrMwO/4jp5Btw3JfOY1oOfnL3LhORhXp9HjTPW0/1HpFZt2eoQmVFtQZV+7a
akDqynbb2qZmfGA4Iixve1xgHXJ6t4rRmNXq8G3XNbpPVJk8iWjjQc/Q79M4gwx4GtrkmG8qgudt
54QqGQxzqRFm+YiyIpF5DozPrdZpYVp+16GWvYh84jeKW8I5Q1QnX9w4vnxUrh1jo7iPZZoYwaa8
XNBEYFLi/8TGTfxVFUqVBYB0C1lrK9G9Dh1KvPiDVR9uyjW0LTX7zgMjmA/cCxJez4HwGtqATXYD
5sHKzIbwHcrN2v4qdcx1zUcUNTkD5bgpuyoAsPt5f450v4ol/eersjFPkPM+V+gdiVU/nAgFmtnc
apHoH9pIj42pZQGAEPipmW0Y8Y1olPfmzRx955FVz30mhp077JxtKtgaZu9XlHMJWpP+R606WA9T
Fl86R7qfAGls/vgnVgUhzyFZ1oyy+8uFQpG7gwgIe4pCQ5diH63mRv7u4NayFEM8dVYltl6SlLUO
JDhd+QKWesmeabVGjk8ZGiqroQMSSerlQhXZhY4IsfU6yeqrEIoSdJ1rqsDexZwnHDnkQCvhGhiS
dV/Z8hTvCJKjiWXnHX7BRsLSw3IzMrNYkIDs4yM46/s8pxdwuA/XNhqwVozt64rAjHiDSP+4rNpG
AdmfEHjqZfuN1JxHknLh6I42TpN9QWP207pUG+Gi0t2Q9Kr9miStatBnKEt65Xc0AOD5mvVweNPn
ryLm2R/mkyTqry0uhgO096vu57gTZgJUoN75rMzNLh3Ttv5hlbdM8evlfmEDzxL/TD+rTXAnj7zS
suLxLrsm85rd7uJG9E+taOSuwC8GMYYPZSTN9tdb5R8BX+0IhdaFwhtS5JEsKNuOXIEPCQKjY8+G
CssJcWIjljqQjAMuO5/RRLn3kzSlqt76+kSRQmJ6xNUq5XgKtlazG2+ZZVWWZ6/kp6klrMf38fL3
359BCutwj+A5D+DGi5zX6ie2QoO5gTSttIcS7Os2UYwNxzWLt6cWgDkjZRfugU0RJQx72SXJVG30
hMP/eqmd8zdESaPqRfIzvHP4W3hEnHGWxQT5BpLbFegiMcWexaqqgHngs0fXO6oOFcNFq1wHyjs6
nx6nows+HnsPQ7+2GiHVXm9Zzm+TTIpwKcG7mBScADY0681cJwKAKundfxBczPCT3BJXkkGw9d93
vnlmDScHkEtfKUSb7r6xfm/Agj6vV+uTNc2853U9n2lEeIbjHL9UG3Y33TAj9gVEuX7+n+cyqUh+
HqYqxl3X5OOkrtm1ovDobq6bwpo/Uo36Ur6TWZ9xRCBZ9GCFDj50eDQcA2dTHSB8AVqYIHcSqthe
plaVCjY6CX0r5CqTc9ji3kbXmTmRgrMQkh5qhKBVFhWDuok5iGV5Xf0YeBAygQlZkfZmJSY7Cp3c
P2yG0VogAmPdVS9Uoq9j6vm1E8/q784wqanwJeujJ6O/T6qP+8TGsFKga2qQJZNhQKqtnLbSsjFI
MZ5Jf7FKLgrfSrnrxbH4iZXnRFGeBnPBdlaUGo8xkEtgynM0D1CHC0J+N3Ofuzq933Skx1FnREL9
R382CRJma6STJ79XvKKzWTPCr+87VLkZIs7eqPq4UrtpsxgZ7wAola23ml+6Jml17oQ0ohOdWtUv
qs5O0LWye8r4HXfv7cqmLE1GDrCyosGbPkhJtHcTn57A3VMZcG33DZwNNE7zKFYJzPDEey4d/lpQ
NbEhetYg9xB8Ehx4rH9wLy7KMJwzJ+w6n8r1WY4+LNmozbIhf9XmEG1a/Kf5NVCJeKwXdJnLcSTg
INLoBGuBFv/NRcUryiDMwk/R1BpHKqRE7XZIzIotD9B0mqN+QMke4inEbFC7SOyQwpAT3nk8u9il
0iZWXEXItKxcpkPSqLLAOHwRkCoh1Z5yf4ASXGTFhU3XN4LxkqdlAlr4fQb97fyRhjlogfgtU038
CCtRiI5q0CDCdPKGUJ+y1moJuxRRg5xCNNtZOBrWchc0pc4bT5Now691C1cMwUvaLwGPSfbT7V46
LI72dgCzLj3F/+sIhSorROykXK2DKj2XaerOkdNJG8bEuLgYppq6yFUjgvkdvf90ONUHfahthUpy
2AENRWHpacK+Fdy+3ZD0VP5v2JqalSc4NQfcOHNjbHQuiQAueCzvxDC15+9NqBdO8U3xrXUjQor7
2WSvJpn6jLz9ogR/Q1Y3efH9VAXJxaeUEXdlGyGXuTut/fY5FqfZSTVzjnNURZ7F7lNAuO+4TQHl
0VVLPa0FqXJfAhRu+TBcPOwkHBx7wluHKwCidk7sakW6y6ZnZSqr3HUEcEwerdxbZjA/DqYWY04L
MvogNUQzy4lqaCuxqUEflNRSIufbNraKuPHqJ53aN/Uv4Bzvu7rQZMU/BB6EM/IzV9SDEr5j51Cv
iQv/12g3gmbJFdojrXQpoXNn8wxWuBqUeonxv47ied1KOYGHJ/JmbUSvt08azcs4/s461Ea22AqT
eHTcX0fetYroKAVkgwYxIqEKZNgqeOxltOx8nH5Ouxsu0FtUpifKE5IpT8ahJczybu898+mhH/Qf
BJfyIB70nRsWH7FDh1gJQkYX+5+HyCZJt+lbKz1A/GWwScDexRAzzuTobROovpguCeZRgL/MvydQ
kFQLz4sgGL6ApfqB4Eb+YmlZ/BWZeyK8RThblPxBz00MqZKUoUu28/ACZ+MY059uUAVpyBQnR8u5
XXMNDT27Z+svjfyRpondB5/IZMpswiQj7GXjXfhMlOUYLPVvPbSTs2mI8ZfA039sg/so9Xrw02jP
S6xuR4iHkJwWxnYcKXbJeBuZ3JCCNnptc/+SB68dkVG/dVG97lL6dBbdliyjFCabm8uXfMfZHnbI
kXeVZAN3rJqH6CV+B5njAYeww1sjs6XZmntRBApGAozbhKKDymzxbxEcTG5dRnLz86s3Gwko2tmX
mE8nCilAaocUvDquv8Zo7LqBTJxrIS9Oa86eYEAGC97K5wDqKd0WsdoLOim4MJyw2xacxYIMe+yu
+wrRI7yOzlXbao2m+QrjdhVgfVYcFE/q0JD8iHuhpjDdk+clQXspQ6CAXLbtd15ydvmAgMSiEt06
3yILr0LSpuotCHojBvRkrtCWafDlaXvPDea6Hs4/Ujo5QmYtbtNNFFF9kR/ByLunXWCl2HTG/umO
Dv6YVErX+HrROrnyIyoPzruHcX5K1o1sKaFVYYu3c5cM58iKhHr1EADjEuWKchdo6jD9aahsbugM
KFdyDA9t2cblFUh3Ye/JbvBQeEg/yxBE5EsPbDybPvtN1D3UBV6m7EhwVPWD1D7sk3JTI//ljMMa
t/eIJH/AURa3/1RN13KNRTA+BiAyWyfcH77XJpiooOtVfKQfoCp7EJziKkdQTnG4PmK6TINYUohP
XZZpFyHnqIkqQ9vUoPGhx+NPxIY5PjbH19MzKC/s79ohurS7C29cuJMAOrCsECVU/EiMSWgyKNB6
WVOKVjXuQ1ElGtq/xCQlIbwbsyt62DBcYENYBxdTCZoOHBHCk871j7jYYRzstZ2oGr+cYlzx5cQx
gCCYYNI3O0Akw6DLTLzpafS+1wAdi6YmZh0eyHLMJtcybNQ3RbubtIIv2Hmtn13ZIEB5oAh2hU3Y
o2IRy03K0fxRxmA0D9YtObk3Eu7ffSZQak6vTRa9Zbj9fkCjY7LQPjD+ntmnGQKd9S+m7ybArdCO
SmHiePyqmWyiFHsAkzIDwRa/0XTFeb13Fs0WoOVgM0Jkm2nM//ZZBEW0f9/YJF8Q7F//0gYY3FfF
pJa5Mc8sRKdHLyH8t/b33B6zkt6Rnj/jxaTE23gtv9EYCz7/1uXu6WNsgx2AWMt9XJoyi/bmPyIm
DqRxWBAnmYhGL3Z1GnRF51N9b01wsCX32ZXwtWDlMpXvrYBbHoHcJOJ4H+A1EEaQEWCDPl1V6zCh
WavnYjRYbIMxrioEi5qGTcAlf/Y7puqCi9nnV7UL0GKLqV2Bhg8o4Ji5MHPrdTJJQIkiXK1SHqHv
xkHuVofvKpmYM3HzGqBfoyydHeXdG5G+1mjztf3x6PgqQZklouWAZ5APyO3UBktwMBPXABTAptGr
nb2fWCKoIP5iJX69noTTt6AyiqyukIAxnDq+OWyAF3PmsIBBFsSyziuotfWzJfg1Kn7MLBhM3rG0
JAlRFl2G5PkmsPMFNlp1ui5gjlkvuWbp9/fJqFkM1wY36xtJHGPnkXQpTSEzz2gW2EbocahwdxFo
YAHXjyH6Dq51NsnapOcoWhaIG/6C9Zz/w7pmI/siIe7K06RcTOHzNBvaVcoavx6KSAd4U6c2S4rz
gbMYCHr9feTjasOda/bdZQFrrqjV3YJBNZzvpZgpKuWhivtasG3aL8hfQDOB+ROOLvmkLAiulX8z
S61a3hmtl7mrCgXepLwidLFsM3iQEyUI9KkdvW9UXwuuCFS/kNHL6I0KqscKIdE8L9JbVKXvOOaU
I4jUzfZVFtgZOOktaJXlRDT4sDGAbWuMZ2hK4c12TKu8Nm+goaqiIr8xzu0cvl070ZL4DoJ3dmHa
kB2TFas2yIBEvGQ9kIZZhC6vob54QtQkXLZg7okE1QgvIrL3IOWhKV20YI2dqEp3dGggkMU7jZJZ
6lY9gKJG5Im9HGB9ET9cCFsCdTATQi0CUXut3FcMCCe8TtD/vcUXxIfGhOIW8KotYcR2lNuWtM6r
e9Yf0EQiutI5leKSEz6Lp7KkEOvU1KeQbkmIlNt6hc7bLdlJD9iUy9It7Qu+2eFPq4RiQsw44F8F
AV6Pz/Wepdb7TYG/BGWbo/js8HU9f7MeVMVRgAUcLY4C7oLE5EBwSkn7M1zcUBP67ZzxrHKRehvH
ZaFkD4cYZpaLwJd8UiX+HcWSLc1BkryY6GsHPMAzwgCtpULS4D5oVT/5EuHnSXLCN4IBDFbpLWz/
05HQe+hgk13Ro6uyXH7jzh6COf5uT6wUKqWw3wPBEn8elNzAbxyeUwX0Cm0Ji2cHTKh5TgIOujMA
Y+uKnDbU0QVaKQlTMVNBr2nh1TnWEKCzY+DHWwzhf4K1CdPwDdSFaEbhHJikuvxUzSb+Bh1Mhe5o
QiN1MnPUj5oTQ1uIOwJQnusnpVRyHdIgSeB+2yV52Yi3S0/XUXoT1DBEy0eNOWTSWBjpGjSlswyJ
6ryjEnDn97n1IlUa9w0z+V+Ccxor8UdL6Ux3YGmywVfzSW3S355LXGlJLktzBGN44jEyUnDb3BeJ
2vOk6UCD6/X5sSxcyMUZWtwqBvzJG9KhOOkJWVclI7PbLU4svsAI8rhidqbzlHxliSeuVIpc61Ru
mv46Duq2hOBWA6DIsaFGS2U2OqocrhDcNFRohTL/OesSb06zwOilNgwiymGlXbDd3CqPLA4ySOsQ
kiBPxSvfHx+6jeUxH3LznbIdgJnDfY40rACYr2PkNFrpJl5wzhWAy5HsMMJTM4lT9XrNOvI/2Eid
6+qj9TzaPXwJwfu6FuxBDXh1hdmK/SbsYPC3Z62Zmt3nPiZm92fvTysq0JjhY8XQPS4CptEsaRxP
vfGbR/9xZrRFryzYcKtejuGThtBBKM1ksB3R9g57DG3pkGO9+WaXiCuw+eNj5W6r24BlblCJbiIR
1C0mV1taCLHTAsmfZRV8TbSE2T3KZRkH2GsU4CAhPPOjaxPpZJILJIBp5koSPKfNeuDUn7CC1uX8
WDycpnTxcMM+AyWy8udFE//iGbEJVLhA68x4kCpSC09bA8RrtSPqiyHJtBzVVaGUW+zigE4qLUQ2
AutAWWbfL5+cwXrU6ubJ5IU6h0c22tGqn0p7wb8fLkjKpdp+mhl5CMrszjgzQZawh8Ki75XFN4xS
fcc5XD3/ac8cokz27fQMPdHdVsoP9MYdPUXc8045sj/FfYegEkpMXrNhnH78tgz8f+czW+pgkAiL
UaX4UtZ4wgP3k6rsiZtXFnBy66PflfLWEHQ04/zb8K9z2sWPQbwLD2ZK2NS28o6zdCx1OLgpGICv
GRGdsZqf3T6ymFxdP0WCtL1gB05hr8JsFE9n2ESE/5VY0X4h7btF1COr9yHXwUvBWN8aKq2c5d1w
qm4GJpVcTveNGs29hYCtYux6foQtGLGqlkKJkEiramXMzdFWzF9JfAC6RGpp/qoKYrCKVC7Mun+8
G+3/AWOTp/liFxvB2orxB/DlddCtWpjk/kGJtx9wjK+LIXYHK/fjQySWCuZfqbkg869M0rLfgVN1
56d9iogT3uI8XEuFD69e54GezF7Hp3d9YaZQHbw4qtkBNDUR3eimm0up+kp0ML2UdQr2IrwLQ3El
g0XFzUhtUDD85qLlEONgSpiCxSthIUMTxMjOgNE8POd0AolAbNUFn5pPUJkGea6Lao0awfkJKqSt
cmFIJAm3YvsjgMxsXOS8qc8aVh7CDEI2Fh7yA2BlsKD+Bvfk5Hc6fWY+OfTfmKpXYG+GpzY9oiDw
BtqDEUtHQUVh5fcmrWJkJH1MVVpzUy3k01aSI7WZSSAwD/Z0LT5dhoMEG4NU4vvOaaZ2M1+y0xTM
dPt6r4UljhOsr5JL8uSkQoMdmvb8n869E4cL1KIv4+eWJAt6JSmDIiZNdVvGL4Bb0GCkhsdh80/c
R6k+7AH4/sEtLwBkAm4CgFhLHo2wGTxcDnKVtY5X5p56/H8F5LAkrFB2c6XAzbCyB2hcb/kiIktt
rJeENDaZarKzgT7ag9A+vrHLkbo1/6DXcgcbRHGSOyOm2oYUpg5OT+U6MfttjrgMd/tlU0pnOXAj
EXZBp4a80yY14g+EgTlEwhpByan2P2xsXIarUlOkgZOqrOce1QizlURE0vDcBcRG55P4Q3UhK353
z5GcnrX3we5hwhmqNpC6XuYPJN5NJ37o+cJcNsa8VBdyl3dGwvJWL90z55klN8BtvG5RtCHv9bYK
VJ1/QZt5DapygHmLJmXFQOrkPAXOQQopjz2LaqY7GnpU5VXU2aXd553DKwyQKKx+46HT1Wn4aN0l
AwMil/LfEJwfg6rFH3OVqDnyoJbD/NpOw/xqEgvciG8ww2cf/IyZf5umX9HkSRcXPTkbDGPARWXz
i/zcPuLq1+FSQKhspujik+c9w9onZkEn0hYTEVPfIfGFUcNTzY8fYdkeHxUpZXfyYprotlPN/R37
zEGYvxzRvgjLdai5QwnlOu6WxxmFPhg6C81O0YwhB/nu4lcgT/E1+Rv397MqJEiwN7oV1KG33pR8
vN0RV2va9JX5NllKV+uBqkyAlI57+FZwhwmA2X5aoIHi1QvJoGvK4iUsMZUKAx53rB7ouBkIVXZp
aBmYDvkuVcZrcR91QPTQxdY4ln5YdYcO+qbcXyCV3FbN0fV9i1kz07ltwLAywHslqgT3A/X5VFz5
3OxswQ3pCqMfl6DS9tqW9CqzbWMzYP15nbhBmhjvUrfm44tkrIYj6rW70JCKLCLpj1jlttN/HwL3
WQR24egCfvoN5TO8GaeC/F37QaOW5VxnizcEizgHmku7QZkc2HwYE9VtQCQ7bFyyBWsonT1e4cHV
K6WuZUG+kwdR6JxtKhHxPVAZfJ1rkm9v0vh0cY1Q5W5rU10A2PZ1cXVfmsjxXPT7RZansPIA0nm5
MfrUIFh0Qw3DLJg89ZypyE2OPUAYB93WILAXoZiR7S+QkvOWykNvqqvUu9e5Q7HRdqydcONKiZ7M
NMp9FNlu0OqYZIAJpPL2M3/jGAc8IH8vfY5ypujQK3VsTVdRNUb8WIcGxBj0H5bCyLPgYXaJtAm8
Bn4icw+Xg01hRmD5kkt+y/kJR8MWksx7+Mtz9FqakdHh8MkIFVGdgfAZCWW7dlmqCKMA8IeiBq6B
mAQNQ3oO+mAZP0pKPIMHpgkP1J2IjxSWEkz03Lb7ERHOJJRjtLYcO7QpNSxPGKb2OyG8VEZtdcx5
voXVYOklHG+QihXsCU7UBGC8oRB6wy3oJcqoo59cCEEO2oxmDPh1D0m0MfH3Wp/GwDAqIPiRyC4o
pjJ3hd22qQC4ESPrquEBpHzAHUmU89Vt+zlcSiNRF5dYetLYBB9B6UD04e6AFfc82Udsqk1EQBza
A5dJamPRBGloVTF1m4jp2TsMbUL5JWvVxbbpnF9DyRu+gY5Hz8sDz10vugM+1/+bfiTNkc216wZU
pDgu2Wk5Ea5OMIqvb2wuQfMzE0KUbAeEEsV40cOJybsxzA06DPvqeRJOzFh03EKk9QvmQz4wJuEh
AzoKU/Q7KF3NSoV54VYTfgbVrPNOsMaU3aNCxt+otGQnDqoYgTs75X6PxQLrnuNdryj8VvT45A1t
tFoxc1YWOiOf+s/UPt6DdLZhrjUj9uu+nMZX8xFQYMxeT8v9KzqS9hROmV8PgJdm6C4VvzSX5eud
f+uxxD3rqpSdygC2awD1zH+F0nNZClMsblJtEZXihKps7wtWmP9wPMOJc5vY8wQqLACwistbBmNZ
rvNJVT/7yg2BPH5n/y5msGOXSjZyG/YQwTvjE82xXqthaOul+vNpv67/fLz3XWiw1PQvKlL9LZsc
yny3y3OaoW/0UG8laa1ThV2oswEbFr7YMBeDrEWz9jxE8Oi+GgAXJVZ4tEpThV+r0j8cDr+O9npD
YYDVjsTR6iJEGM+ltqqNvO6ePRbEO60PM5I7IZfoaiwGSLYUQF0ELqnWBQFsApTloIXweaawZPes
3HHSghN+c4waa+E/WcfoUVrvDuw0Leq0Zfb6Waxgjx5r5GGAWW/GvHAOhVYV5KENF2YnlTASR4PT
isvVwGlhjkMcpj5W8Ve09RAjl805CVzF8kVARzBBkEmkhMphw0XhEEo4Sj4jGSiOHSa4rLkLJwg+
3cTMwk8f/WJpvPxhq8uU7NpeV3ZcE5mB5aRz8vzJrd+pLONbM30UUhWfseZBMioDJnQahndSz0kC
nSF00+My388QucgQL9pQn0dos2za2t+usOykUu9d3q4RKRHQUO6NSheV7mluXdLjTbeKfpg9mfcS
c5rkNqtkmsDCm2fH2TGOJajrqjBbE20lSWcktolC+rnOCc/IvW4shlV8YYva08s7pUHEmSWFxYtf
Of3/lOzaCuHwlp+hMGumPYMsCSgUUyJ++jQSlzV1efqH1thSNlnq6hiOP13lIkx6qFsninIh2odh
9j9SjV7YEoYAeWdvnuOKY2/eF092lxIMe0jHHXv2Cyn5fNQnaVSX/gLr1cwVR6ZRF8OHikSmP+rZ
6O6XkiC3dlW2+/QOEiQ325xYK4d3h+qGGnbIWKWSRHgfZvXVVPzOERK6sYvNh2zbar3rL/4MzOOj
0pMPYttBnDmXZJfRV3/zyF3ywT9oUWFCFfHcQAtqNaybV5ViUUTLR9LApQAiwY19T4uuk90I1Pox
nm+wqENmgiKD+6OD546iSUhHRmY7Mp18BooHVsoO39uEXF6hF4uyr+6vzZMheOvbBlH22K3ai/5U
0rwwcxV1RIfvfIIW/eQb8ax+0mNvL1WY3bL8m3AK91VTsZBVkSfpxCUlnfJQV/JlxR8dASxDmV21
0Tex/JXTqP9oID2AfR13bE5GErui4zgUjD46/B5zI9CGnRhZR+HPLkMVfpw1GOAAI2JriqNxW2cR
Rh+0SrjN0aVuCNbZQSqhmISZmS0eZhbwRH5YCWYCSTkk3udIlCKq8pNvko6e6vJKdRPSal7lflvk
orKEBwbwi2ToUPQyPELfthwiHwJ4Y7bMk+w7pPkrmuSTKgjMCc/KsF07h2Lj+B82V0TNZDieLpS5
gJAWUdSQlArvnqsoBo3+mtROe8xO/fyZqMaGyU+io9aWD63J61pDEdz5frLxXROvMx5h3Mv1XAYM
xXxhhxhbGkXyPjfFeDZfNZEWRthaErqxEptsmB6ATqrD2EaW511zLctdtTGmywlYAFiYnykJmjzo
E/nTn40FGTezDG7gIuo0R4n9bZziYMHEkB80hM1244yGcIBvAlTy7GNcjEtDbFU9mU3JX50U67gA
/KmVqNrvEEMD9VN6xsPrVMbq9YyUkNRaP3TM+N69EW0lPXWOXSg7FTQlKusZxBeYpGRmuYiiGykf
ZJXcXjQsyRO6Tch/0kyeCMoqv9oX4QhzQ57o2GLQbir6Ef15h27ulVxxNDR5shCI6ZWwXdpUcweI
x4E9yCamokOlEMc9ChxTdolTJuY5+Zv528hhtiWjI5IfFjrncR6y37y12k7XEJxLJaPaeGaMnf4W
SYPRVN0wby4NObZM2ZdGu+Z4U1sbeS21RSPnVI+lXpbKZGh0EB8UY+ajflIHjM7/iCbPWalJ8iR7
yOWb8AiAs6s5v028zpMkEqVJ99pOUQLkMdPzyW4qYXeFGoU+AaimOPwnlICvt7DRJgjKRONoe8a7
mAyermRUss6Epmk/FkwPDJ0w8GKk32kSzaeqTYpK3hqVUq0FDu+9PPQ4Bkol2ZeOCD2tphDskYpF
IAzNNFyKKrlL37yYvalZ797TuEXGFWVx+VH9XKR/7CaJpUdw3uroU7tgszQYy8ASdFQFOSjDkHf5
FSGpWG6Q8pCqjZBaHVhngsBn+RkB5Xycalq3Bmq2My/klWVnLRXfsoO+rHamY82O/Xqoxqyz596R
XXEZpbDj4e3V0YkuGczsnsqUMwLnLC5Cy5Gy6h3GitzOvHlRST3vQD7K0r9GUMvHVQyRpKMlwM0e
BhyixxQK38VpUc8Hcg0lPZHnt9q3CIxh9m+QsnpwPXtPyFGJ5nKAem9ksfyAHbl6HFVnO+nA2Sgm
BMbWpEGbhxr2DdVZICbdNrrTaT2Lcb6UPcxnj1QZsfpS5HtJvJngAxQudKYawQBOOKym6vw5ntav
Vx8HLzIF3LtpCKOEIOdZwwkE4hqLsL6RExrUNPHDvtmWXdtLs6p2PpVpcLU7yb+qlBc3TWf7jBIo
NksAtElyqVclucctb8/ya9Ydwa875kdCNzOBwjhb5U5lpVpHWTzl1meWJ+CAw9K5OfQIYvnySt1I
mLaaEtP1R1WR0PqnOIAZm0AqlbJRy1bZWmFrQHzMCTEw+QRksZR5fNxwMRbynB+4BT3tCxaR26vE
SsdXkzFEjJf9sIK4rBdH1TRHGn5BagODlHIBlcWE1mX+FXVZg71U6smQB9KPRStz1saB49K/zLxi
186qkWSf4uuJwxU/w8KLBRDIzFlYUdqUet7aTxPW8C7T8ec8WG0wADWHL/PhTGN+WB21+4u9LgDk
R6Y8ncwnh1YgW8ZntNmJQD+EKgTgpHZwSETNAvoxQENMLD/pMbrP14ooPcGrUBve18GxwRTm99Mg
+HxjR6YmRfWvdecoLyE/UIW9n4V9yuLhYOSIjTmBESvTz6CXIC4u/+LSrgw3q3uOIYEOhD/PDhpv
dHcrFuxKjSrHA0EjdfZrj2R/YEluomiiRt9H3CxaMWLF2X4qk9jSIK8jQvnkC9HG4VgII7R/S3vM
hJMuB6QUqNL19ROD6ZNIaHudL198+fKv+SBXVDljlM7lFwQ9Un4+c6/DlhGPW2A7dm27ufD1rTPN
QoGYkwkfL7eqilgNvUJe+/EpuhfPFKFxbftIeo5igOC2K4eBKOQxmdkYLXmbHt4+wX0cdRtouggs
YKx8CtWJzMpXEdOkeUOUwpq6e75Zioy0eM9fVNXTXvU90Mb981B7gIRGKmgD3WeaiaytALRvObPB
ldSYpIab5WLvGBvaDnewcG8LR4C/x+Sd89E0BHSi0F4UhaNUV5BiULnkUPrleDLrlWPCZfoTli8q
pxew1m0JFVXvuTnFqZS461QksQZoKIWr/i29ElGvXlYfBw1u5imGIceENzZrUPvEjFDblRp6wrLn
U2nxGcX0WST0xeseKdudZQOn8wHixVwF5Kc0U9Fr5uIqGK/DVDaWlATs5njo4T4kmW30wT92qo0W
tmsF7NfNkp/3pXvli+JabBQ6xXosh99y6MjfUK0SDvuaVnT539xs4lCtuaRJNc2EW/WyectxyvSC
5WmLhdbSodVuH16jALbq+vq1W7TavVBEjkuyot6IVDVPVWwYML3ZURtGHIOsI4gk3oCvD2fInDr7
eotuRF4Sbcem/H3U0sitgnw67fkcG7bcCRx68zAPxOYnb3MVQfP1yat0v5doGeBqvoytx3IjeexL
Q1TnjKzzZTsFxOjqpJlz2genCymprMedEloInE+xSwwU/Pqt3GV6Tzo66DYqwZ2w5xpbfUfAQ/YE
cwDiWXWMBiFUIgMgkJTeB8Lbgwk5OWUf7eIyr+jM761MQNvP8axwR0ed813CwiosUzC6iLv8LVig
9BTP0M+kd6rywpUvo+4rdIxzDfBYp2g4GTe92LuF699F2wxW+12OkAK4NFs9rlJbEMlP1weR3s5u
2+v+WPz5KuJ9Kkq5xiueVkATeT5HIoSUhjD9nHVrMxnFUp+PSjIrXkIRDLrt9h/du6AivBLl2FYD
+osJn21pkGNP1VNMxbEj5axLSQnO5pxRfRzV1TJsMal3Cw2MACIlw1fEvAlY6Ktvbn5Z3A/xqC9x
KLpKqWxlfbBxNkdwWhcuvBVgqNjE7c9PfjL1z0EiKNLBU9QshSU/yEuGAT2hzKWJhjD3gLZ3s1zX
D99V70iH7k0olabOi35V14A3IqyGJXk39aEUYTJEsqvgGIEcH7yGOrXrvzLrN3hKfu8c1FPc1BRd
Oq63IMsa0/Og2u5Fjof6/fbwGSOOOKUtLPngCa2EqI2JN69iqvTjvMakbEKG4N1c5oT88Dr9FxEC
QWKB9RWR9pZdE+obYOovA5Vr81+XYkhYvyGyIkgMpQT0qXmRATzy6W+NVacKYiBbtg7wuSTW/qUq
x1g1z3VKYPunrwtY6OC3I4dxmBVNtLVfWtWwoAk/o6vfP9yCXqGQr5fkuJ71FQimFHALGWUo7m4q
u0XboO9guSs7mj4X90StZZFz8JGjFsmmbnCirJt/UDgvHwgu1mRDS4ZEzrmyfxxgxCMB/fq+sW5A
IQBYOlWpGYwQErLuMjkI7XU6pus3Nn6mklVhRhF6vYmLU07VVC2GD+cqTygm77ULtQEwNfxLwksO
gUEhaujEqyLjCH3eMc/pnsPFOmhthI77O8y510n7LDS3lqD4gcTLbACraw1RL3buqhd+n8A6ZoJb
bv7dy0tUewcclHSeyWjwuq8O0DT8B4MrupleH5SPCGqWygEKvzRBYMplKxSRvIQFCwL0sCQrZqHk
wZ3MvxlrXMlXp4JSy2I1O4FiZy2Rb+LHVRwW5EqaJu2c0OS2I5kepxebEZN4qv8VuSxu3VDTf0fS
+weNbZibb+WViW1fS0OVaFH1Gd1p1kFpyVAYsJwkjcnvYSfZ/h76TgR6lpTfbIUQh+BC15Hzo+I6
ElywJHH4UBckqk4hSBfuicNmLOmuMO2OB2AVk0OLwZ49e8mB9WQa5CXwzH3cxAtRsXCsEhboEAPR
Tbil+mkUqd2gRn6AsPyePNTktwSmEHdA0uGp0wjd5JRc8QMgj294vrXDiBpKhtkPh9hHq2BbERF2
gKq21bKMXUBRZ1VrlgGe9JxNC4/BzWoghw15BXgDuIiUs8FNF/ePYisBJQ0blnwLqHTmnv8DcGmW
baxD0q3YveKGJq3sE0x3z+zicG2xAWq+ZBu9kBofhuMCr71DNO50Ku6Hh9pSFb4jAwd5v7KWMcec
3KcOeGRIBiu86bDzT8Mt3K5LJdAUojHL4a0aVslqzhFJHENF3WIXHL9ydx7HDzeX3XOkTJYK0jbD
YCI2KXME8pOJ9hcrBQLRgUexwJMQDCRszCsF4UFyDPIAeps/Lgb4NNu7rCz5WhlpO2+f0T6VMOiO
/Ui0gcHecUZ6AEQzGRUFGAg9zRyxC08IYspFzZBTpchmd6/u8fhZp5PH2yX6MzX7bd02cr/owLEI
pCLmlo9VmfDoxZHm6gniN53MPaqah2343VV2HGMoV/YZ6ixzvAB1PBgBb096b9/UMc9QEXjrm4xk
XujaK5oN4qOAkxUovklYG3uqRRGpbqHBs212H1jxtV0/U1l7PHpT6pubHG0bTq3vTC9oJ2zIhrco
HghnaaOeUiy69gOigmKm5mmPUdv8vQBXzJ2GcZiBp/lr6bDyv8pAisVUCGanCH241M41TSAFWMEk
G4DpeIxJlCHKOTq55JkcZWzltAk8dL01Ua1qfsj/xvV68tPjaI1sVFqWSQeWFJpCKMqBJNH0waFz
jP8diQ0rF2bOQ1KpaIwIAvZTe2OipRlHiSF1ZDhHHQetjJCu3pWEOQbqdFZAdBzaGY+MbI+1aSu3
PanpCd52iipYl36G2MG3CFE9OmKkQohbPJshmG8nKwRFkTo9U3N6e3QfIrIbxVyMw0g8hKEBhcZp
62iG5uOea0+45Wr402XHGmXTURSEkCttuKXRdhMLFQ/v1+3cpqyZTkb+4Bq7Je18Ny99IKXXA3oD
0ux+bIbUFaOvAuVcX422jFVCkDfVF3jOgKVqP1FNpkgohpHLjLhrFfuVtI8z1t/+XKd0o+3f6iwO
GeFYYuDPwDMSpWS3Y05W39VO/ki1O2sG7LUdKhSuhetYBYD5hlZeoZnEUfecSWBrBK3/UH+aX9C8
BY0VRnT5VF5uzzvawu36vjeT88EFIZqCj1hLQ2K4SfaBQIllDT6PonSEKISwe7yHEO6JOtXr2KO3
dZd9ZjEicyBNsxK/1u307tmcMiVVVemAen5/hBW28YRjXxA801kxO3PPIredOv5CYFIhAxbvHj0s
2/uG4OC/nPQDrZXOCwUohgImTvhNbWnq2vLq+3O5sgcgXamD2wx0asNYoi9ZHcj/DoegpNz0lh9A
QZ4YzLPzIH/dWXLQHXK/9mmRv4NpwpB5OSaG4BHULRJq/uRhPNBq6HjZ5EUKfhkWRVmc8JTjxo7J
nQzJRkFqrL1eEo1Xo9lnUsxDDY2W/Y6WQXE+sWBBpBiFtYiIDNwb/M2NxPYlcNVuUPulk3mQ7jBR
Hj57y5MuNa9dsIru7/GBq6RkepdHJ3/4cYbu+HZbA4/Wz8wDuU0uPwRfn90naH/ytxcLVy5nHNLI
7Bw7SK72XQ2Bj4BRk6h7NJA39DNfjimTpOBrb87Nizvwg78ng48Ju1qA1c/ZLmVvKrgCvWimrDJM
YkNp9nunFnKQulMvBUP58hkje0/cEAG+5ZytXCdO5C2YW1fkYRo3EhGtenwTJj9zuIah4zTBD17u
j43g7hMygkJtFsTL3cEAADBaKIinIJp///2tHQpDMbFOI1TAKdMs5yQ9k5DNSBFgOF5iIKB4H59G
SzXsZ6G4V61b+1NYR66AO45Vk3aTEXG889IC9cgV5euqH3Y6ltxRCyIECOIhp4jcetMxj7ErXrNQ
DPK6mRDP4RYDOiZu5W7oV+GeZSjSkw/k4fF/3h7XZ5guU+RaFjz4dKXBQAym6lBwYHuxFZpNzGii
y55nwEP9ngtY1fgslDier8tcYmfrdJO4gXe2aAzltR+LKsZQtKdeKQlnz+o1lCARixp3Yeqmeas0
ajgmteta0NuJSota8oLQooG/B5AdwKYP72kyXRvNsd/nuVeEX6MfyTmEPGzHBk0XECWYe/e/bgHK
SxoMKNoq3/z+67+Bv7BUXy16Xwy3qkEDny+fkCqUA4v8tFvoVV6FUxjAQ/cujFFyF/xhrwMbnjlv
38TN1zQvO1Z5etPzvJEcswOWgpAMLQJBEZannt8HsKdpm02wA9NyLI0QzKdx0wqJNBC3DRm0OI8u
f9zxtQXYUK5hEhi3FUuKLbGLIcoJNfQyfd9A7V7kPynGaOpcH9GSC/l4MvDl5QJ93Qz8ewm1eNde
q+E+irAhPlCG1V2Yxp+/VqdVP4TzoBvQ5WXliVQO65FuFPOcGTeX6BgahSKucUoicGICK8UgsXub
HqD1nqpcsLy6VkywDkPDruSuCsITt15NL9HI8iIgVGtgAnG64tKBC5BciUwCKi7xSEnTwsV5oCMV
BZpyAjIcCyfSJUCE7sOh2vQ4ggGL1PojfPLE+ysf+lIpuRiqekONpaeXvuIJ3ozEgaLCe8yEwCPk
/gkl7WDyM6nCYBQqfhcA5QuPpWr4eHip7AWCQdHtjm22J0dEi7xQP/CQD/B/qB/RP6Gbk4QWzp8P
ORxg1nu9OuXbYYuelC30cBSYtMSjnScDCnE76MNTsO0S1ub6lFdLod2GX1QRl0z19V3mKwTnZvrV
5BXZgRMFVeKsyz9YGQZapAUn3ktOlnbFtXXTeHY1sqNKPOG2FzyYV437zpLlBkqOyhyeda1Qhyr5
VCDvymiZE38xKhh7pzUH42F+vMkJjyDG+SGO41AQ10llQ95gz0di+JeCdfvluf3Nlm7hGyF+8Hv9
SuRc43U/WVJGXs1SFVHL2TlUn4oV3XvxRwzQgnqC+/pLBFhPucFNvfApTF0/MqPwXaPAlPrb89mq
jwyMCFzaemM1eb3lTb7qUdd3RHs/lCB9bxFomKD3WMW2vm+roInzfCmV/tBdsvpjwbH/adyOsCoQ
5w6HpisUHzR0xoGEeIeLXJvQR2bQ7JiGX9TJvykPtoTdQF5Zjdip/GDdiTxgPUblmLZoxXpljk58
lobTizMTtdZPOnUtjMTwc7VyTvjhEEpwHFVwc+NDb8XwdY7bncr6sLNwk1UUwi+b/i1PFPDpww1Z
MRtayRwhuXxhLZ1Z6Z4r7VtazLCzj6fZ99qMf3PTesV4Gv/k3yi2EPnuKrxGWaTWrIf1ulzwwvrU
YAvfGo9FRF6l/yEA6Jl7DqS2K9n0tZllE+JTJLH+r5DwiLhRFTXL60n7fsNsECVlOEpO+sYbjHY9
v9gPwWxznnriRzQKpRX2qjtxqFVv+AjzNCUrpwFn7NilhQ8mgxoD6kE3Xq0MTWCB2Ouj+EJ2MLhY
5xH7O07mDIBzOtawlqjOFm3G3py05yvQKYto7Dz0EHilYnCWd1QaNk+bC17Y/NKddw3Sofyg6lYC
BY9xHGyBQ2H/YbLrYTBETC4FsyLxbYp7cd1vNCNXmbvTn213VFuXqbp3mEvItiSNnysXBZOYTr/i
WltiUYF8HWalLXWVL8ocCm+NBhb2cmMObhW6gdvM7acjgtMMmmxmQXJLPneA4fz/EW4LoPTO7JCx
cMhEUYBE3nXHWcLGeaQZsRUCMeoC5xBrJ/R5JPTPrIYdJ7d5t+4jRB2Be01YCgEsEai4c+yWo3fw
pZZgAsymNNr4T+Gfsm4WMyU6fFR/3vDENx9lBvTg2yPpvGoHcqezBqX0tWDGc48KtbFcSBnhCErP
iVuRY3Yb0vrsO9F6yphLKv+eWjqSshkIuxheeQ39sq9SFvElCTstpYJMvQv+OF3z1uffUVaAgkqW
pT0QQGxOrRZpk9C//0F86fsM5bogKX8JVPcK5upDJggQNCdoUu2a/nZcUu5ATAmx/8XDOG7KIHfw
7WYv6I9OEJdMB6w7gIU1IITaKu4JR0YrlI6tppyBbv5d9f6gvMHuA6yc5Q1wmyAauJelXyR81P/q
nXj2FJzWP4tB1opo3lDVWw7Z5lBjuoDd0M52wM+Dx11I1g+omZ4CGpgriPAcJd5jFRBj8JU5bBxu
qi2DFkzEivjCaE/gHNajErUMPRZU1XTHyABcBoSu/FSu5TvnoI6/VP0DkiXtfh1mDfYHKnDMc8M+
6QjghmPwGbos6X9u9yWukvEYev7W7n0oDFR8xhYY4DQvV0bJsLtIRufdoLYFrpLHPGL5+3lE56nl
yTHQAWVYNQkhYvTKqjglGTpKtHeG7eqHBxiz5QAUsKp05xnI+IShwMlUP/NjxUwzqDvB+0m2oDZw
oXj+Wf2N+joF0EJn+tZoCwetGZqUEezFac9Qol6yGcw+Bzlg/JaJXl1bWOo0yzWkf2jyE2vmYTfI
RCtbsULCHpy8WRBEXoAbfqkuJn05RasCtt6DjonVLKj11MbJj3N04XwV+HfV/Vbke2bzMueroMiz
NFT+ktVrS3/uJAbECo47l4P8IQVnQ97FE+LX7nwPuzPfVsrCLN7RFuTdgKOVWUg7jlP/WxDy8RAf
tbjrl92b1ModutA4bZGKw2zS8DHHV0SdbAtePajsdUWSpHLZK1XFlyZdtZlpeF+HQP9nq3yImIMy
RTx1vBjLr3HiRfRFE4/u7SjTWVPBrGK8P/SzDgdSGeLYCRFwXD0O9M544jHeLCnhJGAIbxjS8vR/
6AeXXbP8RDkWVQkZZUJXeBFFSKznIzulw7wuhNqGh7+p4aotvfPuYR3dPxg55Ix2sAc0vaaCa9q4
bWCelqk1wTFYa2Ne6FfSmoUBhWMCYbxdTDmTFWOLvo/0eShC3AgiVhQeh+M+y36NRQ0zmxEKjCMT
4xi19XdDjQJJLhdzkCgjxD53rza6lr95FPnwg9JHcr1btDx6d81Tv2gYzqML92NPVLa7QY/ztdap
KAD16U1jzCBVtGsOraOBxb+MNgxyE74CNcYRcg8XuI8QnAZGNcyW2ko7QFN+AeNx0isTUnh40hVl
91+CJ0UyE1gi1BRMQgDhZIdyzKWd3lh61m874FqyInQ0rZPVZRXtf0wtG+FJGyzfrJJVvNSR1LRL
uXi01yquAjHzUycIChpmDE7Sw8mrOYtpGt6qxeQzPq3SnsxGeTtcXwzxstxYdeliQzo8etquDIU6
8rQMCvthFeqMTLC/tjt9OwH4JSW5NvHKkXX8KsKhm0ojIWOvOJLo6Fd18Vm3PryyyP1KsIYSSflP
ipdhLrUZio0A4//Rtg+ccocF4wjB3yGfd9QtNNGhVmqvfZ2Iga4PKIOhhPxk4I2Ahiartu/oow+8
GZiY2o3nx0zisHZ8S9rkQ870/KROihsr81cxdZ2y+KgX0FxNaMn/RCT3i0r9xoxWlhbT3NgeWTbK
ty/J9HxLE1qaZ7VR3QwvvjA4aSwmMFP9KGQeNLpc6WyO59Gyh2jfbOVxFhEs8A87jKJFe+543olN
yR+GfHkWh70Prscvabomrg3nzwF5SRQA2D3ccMUM5sxTav6ehkwe3Pt60X7/WtoOrQHIjz5f4v23
p5jmIxRTKcyifvrP4uRAUvPprsbA+yztQt/SlI3bMWiZjWLEKuI7iRi9En2MH2eGfiCdJiqHYNY2
OarSA0Q7FyVSk5immwVnF3Nk3U7YaweIW60Ellry3PPcNAJ0GG26aI0d4hef320oyjjPiByMPFTy
kLnfhD5aUF8EgTe20nDp8eP39/T5brRUdcVzG7ivnNu4sNvhLbKJw/ptU+7IXJ06cXyb0dHocsZw
dEpktuJmrpC1/OtbhbgeiEMw+7B9KShnzzj8EOhXgbCGXBlFhmPPupoGuRZlMUAJdJGkFNrgk3Ga
ec0LmfdrDVAT2ghi+WrfB3Ps7LCXZ67sHhq2mBExrEHi+x0QDyFLwOLyGjGFsMBq74g5U0vi7M87
0waWicl09wI3cQk3q7IoYGAbHWypKxGT4DL1WRNCRb0wRYHVKQslTYo/P+aKLT3DddMsINbzAny2
woTdC+GNlAvDG6d9SD2evgL+JxvXTe6KsEAs0Jn2reY8hI37jpWC7D1OwZmbYRvjLKTSSR3mkiS+
SZ3s6snec7jLJA8F2OOoDUiqIDkb6R3XaWOrkfjPFkOHAjUiCM9u0QVIlDSlTVBsrUqECUw2NHp7
vkLwIcrF9Gr8jTZrHUo6d4PzOIUszngogx0IDIu5cVhi+4NMRhKusFpdsX+pQKkUtP4Zy/+sv+nx
rbKDqgmoYaTKtv/WhZYSnlqYvIqtw9yHz4MZw3bdutkpLT1v3tC0NP031DO2dX9T6MQ8Y+FEsh0K
BPTkvyqXBqvKcKzonodiZgG6exnijVp11TefMl3Jkv2PRcESx8EfzERDUBoHVRXIoMTEa9JBSdZP
+LGALHk1WZt7h1U4xF4w8AsfJ4TySLTAM8vagpECh0TXajN1RKPK776M1d8cUSFcoxlAFKkOBDdh
k2uhIeRQsZjLtqdBLsRi78V5DxyCdyvjc/HzobEvc8hDHzeILxLewHi5n5hhIWNJfrURuQM+QSoX
CNqFUsB5Fd2tNiqVGKFS+g/IsH2XLZ7y4V1cKNNoEFhVF1fRO4jVXDtG7UIIdkJvFBKYvFyskXPm
xIhBx1AKLKXwFc8okWA062ZzcW7aiNSepFNls4AJf7o//I/0At6rg9OQijUy1+N7onIQOa2dl8qx
T3FPUY9sRCQyB6Ayyxl+4kAM130PyoVbxKcRWORB7lzQWJqIRw237oZI7S0o5TEA3A80i0Yop7FM
DxEmk9eadsWQmG1DmoHw5dBZxJrcMoOghH3L6XhJM16LL866nTZOBrqgKANkFGszgZvLZhs/FRQ0
JlZLLmnwboVGQicNTSe3qdq7bcTuT125uXqu75Ycc4FblOYbQEtmbmtYSQmq3rwKPHrIL5ZrNl1j
lvc+IDuiRtbA04DZ+RqMBQicFGh9MqS+boEJUinDRbuvr4hxXEMyHzjIQZG1uq5pu3RqFkK0c2w3
69hijddz19GUS1EIkR03KtU7w2MKEjjV2QMVOoqa/w+0u2GDwVlnYNeAknFNAz5wB4MOmnv1V98f
Zu/3v3NpU84FCa4ZyEVnJywnS2CWQDTMACHCjnzLIs/F0qJhR2YNZLrUhmfVCK+BTNVCKTMux79E
Y6wLQyIWePe2UST/asWcxOFqXc76L0WoB+PtdlcdoSnAjqXkZoytxDNpBU4IUYv450tCCqUBiJ+B
hJ1HsOUiYkV8mbZgV6zC5ec4k/JR1OzXj+vEgT8Uat1LNbbicy0dqzKrNWiGrHcayDFlK17FfOcC
xDiJYa88QR61cZXXsIyfo1xKF2TczqckjFstdMjK3WMbfkCdAJVXPGYqzMbFD1UFW0pum6HLqYc4
WuEKyddypUGfgw2bG7z2mCNM+WCHoqmM7mxJwCoYHnh178wDrNjN1XHkq2Osyohf9GJTNv33oxcu
Zcnxi0lqe2ra6fXl2BOjxWb4wyhcGaeK0F7fXNflYQ3p37GGokamtv1+30i04CBUKDTG9JlXoGti
54A0W3Ksb5R5bKF4bb6MLQgk4ErfGbUFBme+epfJ6Rq4rucsa75XznrZjj1qO1PMKnKdTxYe5Pyv
cvossQQxfGEejpB/h7vj2GWN8hblU5FBMzf4oJtDT51PzFGPK/dMISG7Nl/+D8zLXklHVhGXIfed
siXbASjEvW/e4AIkmREEarN8jzf18xfoo6xxTWG6GCZYVPTpLx4WCHBMDVeUOT84YVdqS8GBMNFl
o2GbbaBKOq3EcJiPOZ0zxGwST5BoQ4famSfkpRJXn8rZ8MvHC3vtxpFqaKXqDylk6p63D0MGzs5X
pFIEkj05/VYksKo/KljNO5YgF5spgMaIsIRh7uHIHi1BqMK3e+JLXIXuN/B4KTc7fXU6fRjpkG9L
OlBse1av9sz2USM7lTntM1Nv3JKWe3E5aBZ6Etdwkr7n1w71IxoFE36wamZiG+X0qeLWxXjlqIbF
Cz44JhT4+3KDkrg/7ytIvI1XfBuZCQMRSxKJ87WehPvBxnKQBErXiLk3MeAOWv+7BDyXYzJuaAb7
bSTqZw+qV4F6OHhLXJhsoYoyOAz9GU1N+Z1ZfPKEYEiOfhlv92ZP0xQGRyvWT9FjaK8ekL51NLKs
daYY8bb5Ddn6I8t3li0ncDeShtFbL4B+dbhm2dutKu5DxbV2rFlUidhY63Rioo83oaRchaSUxUiA
HspZoYrm8BVTXqfSl55wDOr2Sp4USPTsxFF6jkoO3v3zuPWDmZFK/it94nRJrHb6ggxgjB0X5+Yk
utx9YDmisZxzo5hleVhU5MzxdOACfN1DXwPYUt6KwzHr+HoABJ3IJQBwy0c9O21DL6G2WlKxCjbz
ZiidO0Q6uVLuxMhEb/p1Md7kAzAkFfQCQ6O+bHrwbmo7cDaP2gQhd8f5pDDIz1RTtP5Do+rO+m0f
9LF1jnFfPdQxGoD+ygbY1m270HqBXc/n3mXUHLX6chlzLWj922work5xJIrJec+ajuGGFy5ZdOQi
E47c6qVwKCbHoTfWm+dl9KVE0OT4iT81Nb2dUikTRKXPdBdDY4NR97RJ/nhIMo1mi/wk8kAElvPw
pGkx66er0iXwXeO/6Xz0Wp+pfTK/ETfcuAeVNHRfvny4nozz8Qpk3rQSHZJNEKuC7oqx6VAGHD40
OujQdL+wRX+acqSCZn4YASxPH2vxhj5Y3J8IzURUOtAuA+V2nt21qe2aY3pdOXKQDOYJgYd3kjfA
7rI0pu2TeWGxYbvHt2vNsFlN8n8SD+Pikqpbo3xBPoeZ25ukodpSZj+KiKuFp07cetSZkdtTMq4E
W4tmXbNKcvy91FrLWvoEDgcz2OZ7B3feLR8/vBvRpBeejTRqkhN412darum6s8YfifWzQUSgaVMJ
erXbnJ49CAToIGTfS3Jfz7doAkRwGSsX3o2xxy5tdQlUeJuNSvTTrpnllu7bTNHgGgZgPf0O3Tav
2K3LDr6m2PPaV153OzYkPke1NJKeDylwEIZVNqJwWTq2PEIXXpgLH/uGKd6jdlEzGuoTcNMs68kY
mv4DbzzBb9bp23hfGiUNVkKlDibIDmg9fSOOkCAfnGAG9GUlZyIxphRKzQCLC74TZiAfAN8xIumZ
QVQoja9zWd0Lp+hdCJrTLdhcPb2iI96IlEI/HO40U8a695zenoTc1d6zs/7KGD5bdTfuWtGeMH+V
ss44VmpyaixQdVmcN5oAzcV6lNgFFwhOZ5u/8jvZKU/3U6BmZMuOHValWFNDzlSnzJOWxaUtJYL9
4iDaglxhFrPcfJppgdneyLUrhuv2aujN1lCkMwFdqTDqZ6J5WLgE4B7OKNHYs3JFZijDj3sQjykE
7hufcoXG1CIFHZIj/CiTX3V8pr7wJ28vreWDmIUNPteuJwyfCbjHkrGqpwnHekAxJsl578x4MZUw
T9Bt4DOyHaHY7KgVT/gCujoX3z3iDd1jVT/VlPzNooWqUoqxDCOcUdlwROl4F//Z2tMJ82iT3Rg5
WyLTW1AvMEf1MNH3u6mIKUQo3+AJR41w2FxLFBmZTIkfwRyP205fOBFu3niRcjTYnWGmr0feyH/C
b9DShabHF/H1zsgOWawDftawArxkmsMa+/jmB483U+0ISABSVUWNH2emG1KDamnn40mWjG05Tjoc
v2FgiAFlR5hSKnxHcC8HmjcO58a/DALXjAio97FaBlagmEaVs/XWYCAHAUkf8Qi5e24qNbKNbzuc
eB5VNzvPcrhpKDMrkk1kOK6tmnHpS6Js8Z7w7TK7PcMVn+/PtkREWVZ4DkFAfOQ+gihDJOKpmSsL
mJLOGtEgn/yycIEIXFBml2T8cFIaw0QTPxgDGsEQQukQLAf74Up+lw3kNAFRaG2tt5vRqcPwZE93
bzAzTQ2129SIrqKbmBC1nG1isJXy426QveBOIT6GDpuus2oMZIdRQ8nZusLHT8sMo0SAqU7i0O3r
U31yZ9jmKg6p7uF6p7CkQISMY8RcprrZphV2qU0c6EiBj66XIC9HzWzpCmKusI9hxTe9JscCxT6W
5D/3C7EB2yrVJOjZulx6nXPUBrRaboJz5NwaFWUYeNIusdpQN4igaq1EXDKzInNyZ1JSpUwexUrD
wu5mmoZku4c6lvQUhyKtc325vVJVswKUh95OvN1IWBo36r80JTtOWNSsFkVLuekZYe9l/IP5mcdM
TDUNBnXdekkypbKzDuBShk62xMCHPpOIiCbkCZPkSVVDhRaJdklCDj7JoIX5kctdTNGthkp+4h+c
Q+fJ3qDwzwahWLGkyHwxw+ogVxPg0djXG+q/l9NbvNYMtqzv9QpM98Om5xgrwMWN9AHAeH8/Y3oX
11WfqvaPzsTdvAq4UtlZAKC2ZPS8SDOjNIjhKLPcOXS/92m7q1EvdlvVkAVMJ3ccbQi/bAhsiEA/
wwBHBTI44GAfqzXNTEISZUy4JwyzKhON4cvmKoZJePOh2G7q4l3o/L7+n+mFvXFDwjtBY5ullwqp
xVktAhQoYPLhuu3N6ybreNYxG8CplZH0dF3EQI2c5dTQtqmpr2LtGTiPfEg3cYw9S22W+PqvPKrT
mXKxHhwZvTjbXQ2KCEGZiLA04d09volNafmDBfvRKX99YZJDAh36I4gq5OhWYOMSBBSfMOqsUydc
At6HfojAM0L+EiX6k9eF+s0ZEpztEzdRZqqPT5TAgYfPeDcBt+dphv/iC2wftTECo67RlNIHQ0AX
euIpFF5tt7TX7QidKRLwcZk/dqKjXW0pjON07f1ySqd5malc6e8N0qBBQXsyrhOYB1QxfAV7ZKNU
QyDUnR04S4JwLym0m0WkwboKR5udFCa6sbgqOG+YIZ4ngTcLI+9hUTUwaa/xbuDmD/JTcwGYjYzM
z34kwwbHS1CL7ZRuuSldqXnvx4re5BYrglSDFaMC/SstKuJgP513suBp4lNire0oFBbLTk12SN+S
PC2RzFAjFHab2zEjFP/qLDw6x0fapXYx1d2ckuzu8twEnH2RAdPnnOkKS++8+qt19p4zZ6dHkzHb
RkpuCQb/r7y6/Zw79H5mR4Rj91xp0uqYs8i6b2+OIp3kG0aBhAqCXE0CEB6oinAOSK/BQhQDrzcP
iOgOM54+hwtW6fEx+Md2D3hRPvCWihBi+fc88ip8DAZx4t2/oMTXWBAZL4d3tz5AhYhbzHeZ3EXV
gbMSIhW1ptCWjKMSRlHDZ6ORMJSM2U0+7J8BmQDxyFElUDjkf6TIdZYTEE6M8wTao14dkQRq2Ei9
UIoJd/YtToc2mW0bSCKiHe3vmuGShKHd64x9zAH1F5usGmjlzhzKLuCWlNoxqtTXY/PJ8Cl4rxGt
rI2mCcci1x0sCdi1Nny8u1hmWQypzu3pRt7KdNjbrl4fF4SJV09ABRo6c8Eg56TE+k+TaKmdmRyg
Vv84/T/QHFEArRg3LOTE9yrlvqnf/uxY3w609fuCySxxWCLKlt5/NO3mW6/nY8pibYRKzimxdAJ2
p8iH2VpvxMUOmUOIOJTN4SOi3ThyQTG78mZOkAu9iBw8Pfv0Zx98+bKlpx49+U8eVaWyS5VIwNET
ONnFSdMaKWhqo4hOpSKtKrknAW6E5RkcqxW7KHME7ObNm3toVCoz0U7YEHgQ/N5BLNPAzPTL+uG4
rxmoMDvw8Nacl8oEMD6PEVVuJmaczlGPgykseXP469skVx87GFSPDwKJLcDgR+1MIzDYMdsT+WRp
02BlJpFTcU9PKMfWjQ0/zA22jnycwwJ0N08I2eYUTuQtFfqVtJaKFVeDrtY8H0JTHUvzEbT6xzI+
eiN/esRW4WqbgeoTb8+wJqu7Hw9pB8IiI7/HcAyUsSotVg666VwUqsQhRF/UmBJ5plcTNqiyT5BR
VVjl+VlzwN4Hg7Q1o58CEppKgcJJHjSN341H/EyGhNJ51mkyro5GhmiroOHbxX5Pgq8CbqCGPD1r
ZabhBFz1h1CJ/oke1mIxR8FK4NN3yZGSosuTyr8GNmMXOZ4zkIZuL7vaPHKnY1qRF0rG7wSeErty
Nqblhsbc5rlUE99oRm1gHguK7d2kyWPMtrHIN+hqpOVfv/ETWIOcdnidZMKTSrb4r4CbcV3bVwID
auLTSLWf6Yf6N8Xm1l3H0g1uv78vSYKaVE+YPERY3NQlsAlls/SDqNS/j/SIwFgh0DJ+G8r1sDKm
+pTjdVtOCH4jh5cG83A0nnZ1Bd4exfpQjA32vaH45MlKaNSiSbRr2hTysq0ZsQT1epWNm04HL6kp
ZC+q68VUDkqczOAwaZ3zhB7oEniruCFfnutk/Jqk/BZpSbdM0i6LCp62rYyJzN9lfIcsW+Fyzgzi
GbKFMJkMYqE30I2oAlw4Zkx5sBLS69NkZAcabKhN837x9pBP+YVl/bBqvuYlFj2zSRCq+W/lbkUS
3qd0udSLhEJwGXlpWjvfcGofhhAKc/GmjjnUmv+7tjBALKLdAqcjhHtQzNS6aeXEMdVc79cF+zHI
hRAsB2dJ9Q1IpZaXoUmvU8cSgchySuZSI20RQ/Tyn9SfgsiRWe1tpFFAfNfhyR5vvqCrJqdu5db7
Nk3i39twX6+qP1Yqo7o2OwQrmdt1DcyfBjrSI7YGntqFyn6TzAbywiMHZYId5Wk3MmonE+TYauZ1
Kol4Y/HiVrCSElAaf3+0QSrVyJGHr4RhegBj6+5a+UHqUWAkGHcOaDeqLv9BI7cldpZqLzBpoBz6
gqE5Xb1IZxYcmS9E2m/+99vWYMDmtb/MAXtn0YxLgf2S9Fcgq2LJkINq2re8g0ZmuUVnQ+RPrOfh
Ioqs/bRIkLR79yUIJB7OeCHYf4aezew2xmHYJfTb8zqU990NXAl+XNl0NYTStNoEE9qSAs3N9SfJ
0pIWOVIACA70aIlVYBpuRDPm4FMXYepRiV4p3u+vw1/626Cpzq2G1h7y2UccLKmT2E+qBnqkl2Xu
7L74BsC5FweaJ0SDHW5Y9ToE7s6qZvkzSPOOFDPt2sW5HC4fzAPGl2WylvvuaZToZCOOB/9+PjDb
zaaY5jiO+7yNXTDa2qNwO7bRMmByWLH1tp8ujr+fa3zBIk/wkkymEW90rhOsBLP1EAz4Fc4FS0ZA
h0CxqVVhRRamQjXS0BQKiy6JcLXCeIp1+1e/iGZhQnOOlWorNGcdB/WDUwIUgCeM4HXzcb/ZSENs
upf5v+o4K5TTL8hCjmJPNoCShw6D3axGK6o2MQNPhe+QBEEPgykpMcQt+BCxCHSQeEA86bdB0OPS
NQztqQfyvvr8e2INRyqmBOtzRjAKOKefNJj+K4tiiAEL5C/YQGNU6q1WlZt5bkHyV08MAuuA/TeQ
LETOPnkr34ga2XC0nVFzKQRfq9JPMyN+A29/jdxpjI40QSxewmwqsCXwHpgfmw9Z7SEo0sv8lA89
/GsO2sC31K7CFCb2xkw0PilJu/Wh3WbXmz3SfyRu7yP5t4a28QWuHE5q698pJCdg763sRXyyUN5D
BW3oKCgCQl6k44n8MRRaR6BBMTdjVjMcPlk4V1nccxSTSJFuCWGKomGT1cxacijy9i2n8wWnCwfY
ReJbXDgh+PfwoI1lMGUPGCA443vmlkDb0737Ki9GZe4dLIpek+agKFtX6nvdf6peRcNvWyQxyiA/
iilSRNT6O/nmc7QCAKTPltFHMWV6+ShBV86FawT9XQabFk2M3egWj2vp6eH2oy8GXGp13H9IdaW5
YuEq9jimpuSLiUQTeyL8vGULHAt9qM00p3FUrDxsoA38SbzgDZ9Z/nBg1FVy/gqhjXqUtVkLAuFK
M1opjNaddb2Kb6PXgwjSp8y21uQ0oY5Y0mSCsab6S+L5gmwCD6No5Dr2Ka51t+OJ2Yx4/JnGoxpl
t464GPbTfnbN2T/iYN/aIMHnZ5xUZc/z7ZIRDlxu36aWfpZ3R6ztyEfuAw41X2N+HtZHy/LpmzoE
6uAjQwcny3gDHG9DIJG0dP19MmaKcnE3706kzAbcg3ijQlCvljhmMmG5YY4+WFXJVX2rka3NH+c9
UsKVKL9floKybNba+h4O6s4SnPJFj+3Slrr5nn4CbMIGHq54euyQFbXD3y/AcRwbz+gPARZOpG9f
Qz1PQguAJ2l0ynsLC8t/KcoIdkEYhgDE3upv5oTeRPlx9aFKwv+jrezIl1UAIeSspveuhEUfTm2n
kpf7KOko5icPGUCbsX3pre7MbG8KiiBANo4Jf50dQC1ZjlsPjUMNPMrhWCLAC0I0Eo2aIc0oOPx6
9yzsJcQQffPgnjFHRRxJ981jjjNfHA2VAzAJhgYkxWFHFyfyo+8bOS7scwZz27JMObBhw7rkOXrn
6SydKFId0woB2L8ylp7NXWAnLmXBTiUmB9I0H0eepgmg1EQiVV4tyyXyamaZ5CQCsFGoeWgxNeo9
Cme/7Ego+e4pHtC3xkTfmbGcjTKmqx3mySYbr2NgqOFh8dwfWkwqA0ojQiYM+YAaiyuz37jlAENh
29awOYPcIvpEsgHmAMzarcgG/oB1TZpVstC7jZ/zh9QHt13v0V0L8JDPyJ+kds5z6XItlmJiscOd
A635PO3JXaBO5u2t7ErdVxJ3AVbcMCyTEDTnITLsKP9VjVc/xSt8Y6uNHLRmKjCTDplonHgNVFDt
pgnApv6GP20YtUnS+hNeTLUC2XDCk2iHZW+pjiBYY0Jfy++ifOPBIZgg5llE44oMIu7uaO3o7wu0
QZYWH9ZSOfX+3hoNwGEYqeOi2giiLo6Ve9MMXTBnZQqbeYYI1qQeEaJujSkElBOax4kwpr02FRz5
VoWlq3b1ODsELrNzqNHCbcAUv0RzEY0q+KvnfMVmRlUwV7MwVpeTOrLszSKwNdweDInOVn+Z7OXZ
SyxSrhbQho08T1sm+sTGTCaI1g3/4LVz/1nbP+cC+8goDflkq746qFvrP4TKPWeCqCTRkbiG8RVY
N5GHl2l8kCgSUzlcYhoMWzCpTZ0qq4f6z5LpnX46N36M+ioYqlYr7mX42nZm+nX9mFpftFvblfnu
0FDEV1yv/cg2KiFp2F1cDH3RIFtQb7ygYuJzscqrPnaPEL0x269TiNpheq5LbROKLM6uZGrHeBN2
KKBZT2WEITY1V3z79nE7ZThcZAoYlTel+5wCuz/WK4MhtDyyhMnBUA+PmV09VKsM9I0h2GmjJxNj
3QQOXW/0PTcpOQfxf1rq9IsRZx7viFOwqpuVAJpC9Uwt0MkCz5jA4AToUTDIY+igb9fzwgzHpPnn
dLV84uTJz473ct34fwhmbye3Ej9CgQiX8lNgVxYZzbsTFjxnJW3j4WcSlp9r90AgYQQB6NEGjOxC
nVjDPiXcyNvmJnl/8cztPG1ys5bIi64j5V0W+ZdvKrRx+6SZJbh/S+/WpaE6veW1DkvLQ/nwYBrN
Xan+RQoajp83S67HEXdO9bFof16nM3CsWQiO9uOcv0ldZ1eusqR3oNk8SmfpDgeyvZXGXSWCLWxa
ljCXAoIM6S68C7prfHl4ag4TwFsR9LksHMYmu+HwpEd9TCU1l0G9QjitvWHqQyJgEZcXaoQf0CS0
lw4iTczAAkQ6a+Jjmz3PKFMcDge5VSzajy74JTQhHANm6q0KQRLg5G1J/WBkIYffnEkl/04fg6DP
GczCO0jf7X6AFRYWYUGLJh5mox7NqeSByllqhJJ8nO56lzm+Fg7O6rZxb30xCGyybJXVQ6whCB7D
6HrX43MwX9hUAtxwaf2S18QZqTrZNWP6JmhiJMST+GIww1rmKTNI6n7Vk0TCZw3X+vp/HyivyKGH
WAd/IFa92pdpjajDKxLcZcdHQUJQJsF/EcDXV++ieCgwlAcMkZsR97liuIrCB02M2s6EF1R5s0vt
5Quo8UeOzG4PVnNtWMWv1R9nO1skzvlWs78/ykeRDe8+PNhApTlJPToNsjRBzMLRXv9A8fswaZR7
TrS1AzeSLdi85oXd0WnqvNY9rkuG/R6W9nJkfq2bvrFnpWAxJ7FgmMOkAmfbxStrpbhdORFdkxcY
m4vjJZ+hJmu7l7KyXM+YV84lWTomhSowwvY9B6uacsvcirfG3er1/JjeFB1zY2WBqIibuQWtTJQ2
RcobakGU5f5vdkksn9lVViQ08Sh0dpUk7rh/cBu+6dfPbyFF7Zt+z8fKwCKLArn9ginYUSGgpisU
p0IrkwFwHUCDfwQGna8eS2d83VMy9kluwtExSfpKoi7weiQEMSKXfwVCkuyAvUmbiPTVIxF1AcR0
dabs2i3l7Kr/voBZplZdWlEv/M/BcNeDsAqmQLnRYZlZ/tDD3BjOUED9MHEZfU9pFUnqUE96YSjD
2sKP+gihaHwJy5SbBrq2SJoa5Th8HoBRFxTQcuJQCtzkBQR3llCqpq8a9bbCwZ7GPoEhdPJIPiUy
2XkI8/eqFNgmujMvwzunsx4jMLJ8FCiTEJ1MDeyT18appe9MeKOsGmuzxGd+AoUqcaimwBh9u4Wd
o1PrOj2gh9BovG8FDalNNYWf4awbv8bcCfSG8SiqLjeQx9eIhwZgdXh1e5ncfDzmfw7fzn53vR+Z
XMyBsP9AgpjhGazsLFoRol+HcebgJP9AKMgK4JZRTAxz+b/jKrDb0s3Z8cbd+v5a3mb33NoP7aLb
ZgGbEH6TVMn/7RDQP1pmhyNu1wupBa4ewIP/9E2ZO5Vt+ActH3FiOpNFiR4LZw87N9s3W0cxFhd+
ekIduHnMZGXLY86BcwMB8Drgj3RHmr2Jy/9n/pypmGKrphnV35Excp4KLIAvp3auLnU77Y9trra2
yL3yjmeTfrMeeY3TxHvKolZzfq/kTtVT5Cdfn1j708UFYCC9VG4TNfQbHKb5MrRelbVG2nwxRPpQ
oKJRS54IbROns7R3aeq3iB6ua5bXD6Yy9YRdFCwMxpBVimdGcLh5jJMH/FkwHeXTxxsPrbeSwpAP
0VckivI8KTZvbXb51NrXZHmnleR2rwSrrWLklboKlfj84TYb4MAkSxK+s1BUh8mV0E8CmE6V6oDv
lnjI2BfF/I+//kOBGvvSsxbgUYUEykaVF5b3+rqghX0A1SP6DH7qWff2nkyYC6PkwIIuiTkmKVC3
EoUxXZbhb6+7D3zU/z3fA4DS0r+BdzmIgEfFCW1xOe/BvoEOpVdTcBNmqc9dbz2XbTdxOLVO67ab
omwdGLUhQkaXKzYncmc6yE7C3TRSG/xpGifj7A/U6Ms6+Ylc/yMY0bJNUHdjxKeL81ebagbhRxQJ
gDhJXxG+YbxoKh8oVssWaAVhiiKt1bT1di2zr/6/Bn7bi1Z/Y5aDqZIqjHeUHnjISCRmkTe2/h8s
11/S3rxOf0iIpaCqBPdQKl3fDQiunjt359l+bv/m9y0wN6M63fY6taiNMPwEWS8O5j+joT+nPtDQ
0hvjgeVL0gsqRKGi+2g9yE9nhqz/7K2gJVrKcfv4baXBaHoBwD0yjwoERjUIljenLth/GpoJ15+0
eQdyzuKkanZzLmHtwj3ATN90CwHFZPSdoJNzvc1nTuOTjnCjPVMsdan5uUocT7aHvzHxbX8CnfLE
/9JMagKQSG2WbeoFlxuBginj/p/uKBs94EjuznSkf1YAqTJWt2kYL+HAOqCNh2X/BjU9aUF4B3hO
NBX0PYhzwWXCEn6/PrzLCpgB2HjjEzDWW3n+1T8C9B+xPMQVaOH+3ZELs/BHmNixph+ewb0mX9Vv
BgdY3mT7nXiLJHBJazI24JUXg9r8x5LhcMAPw0gYhuU2Tlp0E8AluPMQbyavOcXHKF0OnV41flts
LY/vy084GaO93ja/ghy/YANKKPniEOzvfJW5KToVZ233hgLzjZVRx7f4rFJjc7+FY0X1sSgOnT2b
z6vjB13qL/SgYJHYbgvx+Da4vtvmme/p2Gm7melWVpxvSXUw1ZsJh2cYwNWhC1aAaXihwNebFQ+Q
otwHjaiDDS22JAgUwkVwI7zjtuK+uYI3uex2YipJmWq7bEEJHKKBm7uq1+Wp+/43PJkUecdg01Dy
6zbZhxJpjgidvmZo0+owFOzSyQHHFEYrBkRvTbgGYu5Vq1Fxily8tJALeXtkcnDY3oe3ih/Zp/RV
zq9/FrHrfGzBSz0D0oR1HVDa9T0Vret39bSEoN+kEfH5zW/EIt5bdyi8l2d6DWI4aSJLmHDRfknk
Spo9HNY3yenyRlSKFKu2IOM6JdIyNCqn5tgVWzJ1Ty4/y96dSP8jZ5JSoX0itsmbzZzXAlHCwT7g
IoiiZFltrwRM+JJ/HNorgBUd0ArCpOkTbyHT60WGMvfGCL05AiTiM1Qxecat5eCaT0auNl4RlQPq
SrjhwZIKwDVpT4eTs/egBjxLihPrI/siPmP3Arl/D5KuaGoQc2AlxFG2WkPL598JSp/eoIemnKR2
ihOiHU6J6jENa26e6lVGH+i4KfDayMHT308pm/gA/Wgpz7wWUD3QrzJM3XqkHRmZB8Qo+z6T6rGy
HXaSmQN/haSb0cptuMrNaE93Q0thJ70+qvYISxqQGBBd1Ur4McR42mKhfU9aMg8m6PB69UJPYwYq
1A+LGk7EhULIHexMF6OfEzKBLjNtg4r2kVGfm4f3HHhnREpn4DF0uRl+0rGsDReAqrrcune1kcRm
/StGD32Y5x1kQKr3VRh9i3zzXzMvARsPifKf+G6P6JmFzPHuL0WEVqVL0gU3z8Gvh8V6u4WFcREt
JG4WREc3DfwCPwvcrkkFMuI8s21ppCePqBOoamnjrqJ6JLGzTTPSy+czxmKCJ4r6TifAcdEaMwWk
VrtvsMienkI1VPT1LjXaruGPoVsGWPX0L4ZY6a/50r7LcEvfI4Bwmz7N7Ipt/JktocBbuyPDk6ca
Lr0FPSKl5VTEbbxIW3YRxLgMGKl8HDmDmIwEU0H1BiigxxlC9BiToIl1PeObTbkxxjlIX09XC+bx
26v3jGknlT0K8mTcqdx0mu84gpBt6dhGLs4K2mtk3zRzGY8gRe87bKUXKXziX0FKyWi2XoY79cGW
kC5mKLmM3i0aCz7UFW3mmXCH4LKREUV2HfwoLYJNq8ortJS5ecid3+C9vy5cku0wQDzGApRLXUSb
IyGTW319MNF171mN8wil3XbZXI5AEO6ecsNeviVUjvPqm2gQXDtQ4BYvQ9rze3JJwg6OVHCdL2oc
U/TV1qsPzN2UA+lD/zLKNp0240elCt8RE0xrqTKCWbO9rwishaXLr7YSU64yNqKq9rsQMMcjjhr7
23UKogXAqC/3PPyIF7wC66GjHW7qxrNkbQVHDbA3BtPesBue1UxWVBgHMww+eN2v5bRY6I5O7lxP
ZC2zckyaorPNEkn3fDHIMPdpB+ahG+Uqiaaz4SwZUBvGs8WT3SIdqCONndXU5CwBxyHJ4zlL/Aw7
+FsaooudKRCkTt5H+hEtNbsP1PjxicBYWcyKqjkgbp6CRmifBoud6lvKIaoo/QNqfvFnQ5DIr19S
DC8voMNwdJyo+gKDRu/ZD/HS9LoLUChDc4puqraU+m4IHjuibwLI2cs6r5mg/8XgDKE9J9b9B4Dj
ighTBox4jzdrg7nKas1uXUGJMPluW34c9ZiIwoNMsm3cmkPtB7j+L0/pjLjf5aBUyfpubwbxX6vG
Qw9lGFn7WcSJQNa8XHi0aLT+EWfbtyrHD0HWm52fx/Rv7evFRmeBT0VSee4ljR3Aih+DP5uGQSWR
p/2eWsTFlWsY9dwav07Mn7I5maHl/dKvyF42kZyWX7/RFspddgsSROaYCJ0JDdFPSefk5rGm9PtN
0KcWCicFIkp8OuZc/9J8eSQ1yX8q0L0NdShq71EVZMv0rkbcxQoMj8HVNjug5aCBx6qZYZGlR+/U
/B0l2z8PxcKfUeG0RSJgClwisli3FHGZJ3G6Ane0fiRGPdrUpkVZ06QYkFeC9K9Ra3aT1+O2sYx9
w66FjnSPo4WrK5rkjV0zRlBHLVgRdTvlYhWzLoQXmeKZgOg7n6lMRfTQOgtP4PPLbyjprbOKljPb
wo15AUyLCk+GXaUy+8KB09iosXsQzK2xigpen0KePWpaIyiWNDmqwVR87XNdTi2hldAp/EnP1+/a
B90U1L4uMAbVJl5cYtf6FouKHvvk3/0fmKo1H3z+l+OCqAQnkGyKmcBmINH3JzryVBJnYRacWjcS
O/6+MlBBPj8LxIMdxJnUdf4iVAazi4HtDlrU65hrqIe7CW6/nSpwsm4lK1Q6tviweM0t8LlGpE9V
kr/2Yenk4TWp5ks7z4QU8STvDBJFCjUink0/Qm+RiL0ReLOTMG9qothCpi8y9y8OhY9bWJvhNVm3
haCtVlg9x2scoSfyWMPtBh4k76uGktLB4n6MDEuwO20OmHe7I327G4hq2Mzgnn5qfNGVOBM88XKw
JWWTgl5WMlHNURhvMRyvgiQ4R5hvyIa9ao80uKYtQ9bRGiQdTz6zlUnP4vbva3bvYswjaW0HpGr9
0eOr98tqu0pMufmkGPbxtyT8yxC1dDcSpzhJvyI9hoH5nyzhl1Mf8PWMakB0QxDImF/2rgSL4u8g
yWCdjQwYb6qoqaSDn6vqe2U2HD63HN+khl3zlBF5ZHHfDgHTzOP655FQ0FlSCFVFxafU+ONrb4xb
sPOuGWxIyJlsRwzVzF8bEDvh/UIuCfV7Y2AMOY05N2BXoFENMQPtXBqyc/Nr2XtC+WE9MaQFosKQ
3+FXaGGw6P86ko1qzGLXzAtCZOuC0P3IqtMnnKQtWaRSKT4LK5tvYKfm7xitk7rJTz4QYatsf0za
tFX8GAJLZB8H82h4xBgmyP1PCInCn/QxevOBBaUqjy3s6QMduVvvSFvdAotYjNZE3qhS4I3kbyVR
s4jEk70hDJoBQSPswJrUT5eZf1JiwnSeMFyPYhuHH6RWXEq7l/M+XSRjonoM7UgcrnNPhvR3j+Je
iCCHdLq6k2IX5dFaeL3uK8P6D7NkCcIsYbDpAYlae7PFE0D2VWeUa5ChN0IFq5so4Gh/dbsjb9QJ
l9T/NEdx5jPmTRsgyY9x9T7WecG8UrcSV92Nkh1kWFkaNlupZya5ZW/6yP0gRcrqELZQ24jjGE2r
0UCmZRDtjrZZpi7Y+NAtp1I+pD1jh0BIXgSrio1mWOPHAe1rvkUiRAWC5JBZFRC43oFc9gvGKnNM
G/wcNqGxCL0gXDPYiMpHTGNQTr+sia6+dFABaQmU4F/77Q9rm/jifljaxXCo2iCVdnzxclZPX/Pz
x+SMR/YaMmWsKSkhJccUnFEVj3WIKOEqUnNRBSJ4yLPbD5QcjeucK0HsOPoIBjQ15lSpkbrgUW2b
xrbDU9w4aZu1yrjWov6KZDjHrRpGGAshkEfdlF7XcYgZqyr3/FU7Oi+hT58fnCoUD/5ghhEHvs6g
15jO68rsB4VPygvdJpYsI4H5aNo3xZ+ZrOEtjX4w9qsIoWwjStNFLJZsz0w3g7gnKRHFQPZ+sIaN
sX/Nc9XA7LzbKC+QZ2yhKy2XTBaXHV3kOFZvwlvHwKztCPTKckVelvxRyg+yAvNvDEMrELM73GE4
zrVpU/uboR2c7/5kgzfKPEF02DX562Lj9ZN0XnHBQOvN9yM+hws5KtWjLWYzvK/3rkWhT67cfrIt
7TgVnm8oeWQzSUW7PNblqD7L/9hGC8cG7GWEVxw8bNMNcyb3USWfhSZv5E6ggnUY0vspKVavu8sj
9pRojBOIi5bLG+nNdrTfzxWQn4YWtFppfYyTxo8z3LWPx1mz+DHPAgeB3rrpi+2jUbUk+w4mWvj8
K4rtGIR0dwiZ4Y7iEHVcDJNTHRjidgXtb/4YWPs4/d5upkZVIh9RbHJGXudD2px3dv8MOAUfh20Q
gXP6xRyDBNA8xmhx97jpTivSfsN0Eg7pv88eR7wTkKAwtDFov5WbrVhTMugFCr8ENQ0qlSdR1VU9
Qiisw4Ew2b6aeBUDXsDP/W9LxRpFNH1bFQo5uL7z56XhZLQcI2oZT00l9eAe4t+Jli2oFrJE+BwK
KExWLwW9kobC0xZ/l4XgHGzc7/MELNonUzvjE0bZV9SZ5TOypEUAEt5J+hho7pjh594/lFzV5aFr
S3KB7DqGvOqCsazMChP1UUr/WlYgsNH9KcVbGa92SoJee8JK8P8PTfaWEr66GJnOBnB8kP4Mcbfp
QySOTVU6efdW0SVxPSp/KQaxfZU+h7hl9gjSK/5jYJWNaCaD7UTPVr6Ocymjf5Vza7bJNpHNM40Q
mi3+n2LYJBuEIxdWhkooaJ7oOXFdu49Fx4RDfAcA7Wy/y4TdLEfa58ipN9oSTHFLCufaXdo1tPjY
0LZw3ncmgySOhzD9toaqVAs7wGMzCtz0cn2JzNgm8E0OofyN5oCB1dPzKoMeOvK8fcempHFg+Im2
xykRw1PtbU5dy5urKIL3vn+AYzfCjp7B7E4cBheBOB0MXhKmwXI9zmhRtiBircwnYz6MQlEQQymi
I2o7jxV2cp8Xo9T6Z59WRy21PE2VSkT+HgLiw0JDcjdMvHt4avnv/8OnprhRin3OyOE6gsGk+7ab
f3PoDZsytKx/PW/QJJ0dKLIztPgm2H61U70FLrweH57a0rX5JzQcnAsmr4pZzf42lYDj54aUDsgl
ZXnd6EIhnZa9fpD8BYU+ankt4M2T7V66RWZZB5HoOgwqWA2lnv7z7k6ufhqYHRLLOHIHSOp9hsZ4
wuzgrgVGncDDd17sTo5vI+4H8uxLVz+e7cHs1EAOpWdB9ohWcSc7AfvUBawg9zD9HN0kZa0h0HtH
YvxX3J5j7PqhPorzq+0VK3RL8u0hJWGV0jgel4hXwR8hnvGbc7vKMcAfjGF4ow/lUvIAtXTWiVSL
zDsJH/VczmeaM1OT9SCeJ1HaKBXSrPANh/pb+r+d9Tex/b9dOZPFXYVmp4SqYjB3XB1SHj3muhqS
Ka6osVTzzHuUwwXsJefBJTUaUCxL4WBVQRrH2wFn0cAVLKqmBCfvZXA+OW0Uf+BiU1IQYLNtIMQn
gYljVpmmkDMYyAfaJiUYFUSFgEx2UmcYDuU2yeOWKzGsyFM80va8fmdVmvJBHYbwFazgU+G7UJnX
Uzj62EzXuSsztVCot8V83T8W+iT+opscA+WWd0A8GZWT9ru1/oSZpDVsC9//dW5lgkEx39hkc+/d
dQMsRL2xyWWg8mLKTH3G48TinVQmznMEkfyqtdcZLuhsmd8fWuJ7Dro8aw0sP/X77Frvmp7XTDNR
PXql0NsGv4vdFbJ3iBF4CtZ2F4koQfcJ9COssaLbETVlMGhCzATyChX04HT1Mto3VdCEr8Wi8swk
QX/w2nNV9Zek3zMGY669iL1jjJGVCoR64KH8cnfQf1EykWQadNKOOKAZclL3kv4r8YTd/+tXN6N6
2bSkpmLcgylwzIoqzn8Y1k5KGRGC+pB2HTRhcrfArzjwVHbuQ4XuGuqoC8zmmOuXM441Ej2MzHL8
PwPmmSeY8Nc3CC1oK7kNu4uFneUAUuDiUIqTm5rxqrVV0wbLEsMa47PNPZpexa07N0MHHtDiU1Tf
lsZpQTfKjPsN0P9fwRhgodqGM59hpPSlpXsUgLDUh5BsAaI7yLNQk/7g7+/a/OTrDFKYWwwfjVgK
dDX12uaU7REW1mx4KGZlSQAK052pYlicLCnzDyLxXUhQY0I5WAdfBdvDOBx7eXVCOndtfCLLojz4
pLkpg8dS/t2e3RrAIJ2tb3/DKFsylcKiP0aNjp7B//queNJtkDYztTY16K8D9YcmzuvBBEuIBTWo
CbgqpcYTuv+AOSdaKu8A6M9f0WQiW4e16MkxrO404K8EmCIzEnNMTnxHOvf2DDZuZT2M+s2xtQmL
CDeKR5U79oKazsj8DaLlt0duZyP6jbYUr6scr30KxvrY4TuAJBRCXtFKUus7fxWSWu7S60Zv5EeS
0ntfH8e/WAtOycEON1/yYo5ggy0ttn6SOdMuDsmgnolDq2r6jqRBULlE8VlZqRun4HjloPV9OfV4
GGoKOi71B+g2Wm+OzuxuTk6D3DRekIJWHC45kM6udjKKCwP7k/mNMxT1Q6PH8s+EjcGnDsudZSHI
BtrvZGkNtWNoZD5RCBk3ZkrLK+8Mn2Ch5nse0ZxoAUdigeV7R4g1LG4khpU2mtLXuGtiy7/aWkrp
CFiv/k8BTXcnhUIP7PrZyGFdqTJFT9/CaWdxBeqEb/88VAQvpCsG1pAtLt7FTqsApJ4+3i4AejUk
Bl1nOnqV80QH1izqUDcsvupKEDaQtLZNvi0wpBx+7ypIIFTLIYOsygzkOmIgLvr6aAqN/P7u0/Kv
nBU6FNbfZmDOhkTbT73FUYsOVsGd93Ef1F2om8AodK8A3PSw9qbH49qUOxAWYWtVGN5tCSkIDlR7
/6GGDsM94emmdo3x09heH8uT2NLj6lr5UAXiN2Pon2inl2ZmYzgOhoba7ySXCJeKEDZtNRzuIYi0
b71hnCzbHq5T3bxJVFf10EAtLIu0nTJFS/Pg5BATa4jDFls8/r5nMdVOwDN2XuVsV6+G27II0g03
+y+zw913TlrfsaamEqLogEFQWOSijmSsNBGJIwFLZDSUxnu5nlHenMaxvAGRcA5nHw0DpIFdDvSt
8V89anEJ/84X6uWHzeKVnk3KcrK5AB9BQhdvS/VCN4I7jQ5qjCWWg/X/kboSL/fq5x+dO11ioDeO
jVb2MfpT/FX9LYG93yIgYpsY5HdAV0Amz3TrEKlLdwgcNtvx2jneH/BExBx3XQQs5BHW6EEafWag
3kof3rhfG7SfoOcJdi9d4haS89yMSl6as+F6FxJCCkaZUOyEAbUjE6M9g1O5HhlS4nlGN5MQnWLq
EWK4LeUPIo5MG05VonqGkPyy/ccwxJk09rzSNmzVlU9lFhpk8xixX6iUtQfduDDGPMiTC39EMQ/T
Moa9I/g5cmW0mgV4PdjrJMDh8d1ONugo/3V4DUcEglzk4EwINL4mK50sF94DSoSOvSmlOc39IEqR
QzIq13kuOGuaKRVE7pAhzVwi/Qxik0fIqjJ/x3KgT5L4Sc2iLuYrbCiCiN2A2SlDv+2ZgmAXHsoj
oSoyKOLeVzmJDGEQM1J/Ske/QBr7me4/1kjqQc5mk81VwuPwRDRx8BQiBjrqPNNzpbyXP2Rn+wdP
xv3qphYLIeKsHS/uF7Q6QIPSuhOZ96ZHI5R5sdkLw8IWgZ/l/whqUnEVLEVpjLzlHpYf7QtbwhxF
Ulh02FIpAcI+5UJwaYQy7T3PGSIAzK9/ev1+/VlRQ34HxFhaZ7LUHoa37W+sdbNyA0sWPMsrJMaY
WTo7ubO0y6d13iGaqOyCZYww9+Sq2Zu/YFx93kv7/0/kxxJRXYOuVFPSYZVs8Lwp9wptrAyVopg6
fYDn+um65buySC3w499JekehlH/ohqQsEGvHuaK5gDO49bzEobiyJZ+JefKeTI51QOeO3XGRzOqs
DzHgY30RDssgxhukGi1PPem+r5tytog6V3YVXmNFwCp//iB3ahMiWLWe0N4FUh//6fi+MwqW+z1/
r7ijt42mxrb2MMY/+x4KZNjRmOQ6Eogw2lwiAxaqynh3XSk5pN4qypVqb4aZrlx6XHWJpyBipyuU
tDY2NIeah1ektIdPmDC8k7UmlhqcDFg6Xwm3Rja18GhwYlT3td6l+t8YxfKBipUyOiMYego1FJTx
oQfZRSw0OYdIlZ/p4Zzs7VwrAdBSvAMrg/51aqbHI3ST+oay2dX4qL/iKZRKHmezCZaFNvh4xAB1
LPqv5auF9KMFX9UnNWUpxUqGL1WEE4F5I2Jp730cVU4pTdYh4BbikaNkWtkkVicu1CnoMRA9oloS
PwnGyTN6xGC2mUB/NzkUmHcdUMj5tbq7hY0i1Kowxjrl3pDU81tCfwszKkaYWk1ns4v7n1e9zesp
8h9PGse/ryShEGPfa3lz2MS2TEOiaisXHjy/xy0OPocatsQTuECh+IsahchEATmbp8eJq7zwZ5T9
fxcftA81hCpqPOCGjKXZ+PfU5D4541KCNwHxoVl0nYbRIAQCCxVw2SxEZx34cbM5xTwOkkVXcF96
D7qqCJlfA6ZtGLibnUAokjc7/En0m1b3hTYSC2nvAT0smzZgf6YgKS1+htLr05wp5wabGZZkZCXM
r8pjMrLXhkft7tkcQCC1rtD+71JKqeehEWZXT7vnDuZsmi1Svv7qP2xx+o7CpxaiER5CfppumJNq
nGBI9Lx36nMdqUSB30daorQmoYvP4gDY7lsBmUgB8XwLec6dHzTltFsKWScmpKptD4NP4H5x2Vaw
9EJ37oZdpx+RAez3KfSJ6G7UODguWLhmI8eHip6IN3eCL2+x5YNR02jnysa5iImtfg27N+J1CdKg
NzI7dPRlaiuaCuw19+RfbGpSM8IVxwwKxDcgugCAmzvigsnGQvkzFCLcb6ZEGWXlEtzFofFCQBwP
2SfePI+nXqecGPvxttyTil5e4UKagqM5lgtV/QsP5xJIf78thRIMcNK+FeYLBpTxfMwPEAJODTIf
FEodjv936FVoWUqQYe3Zov//bR0Z90kh951yvTRGWM63zDzXQTNUb7Cb6y2IQ+1Ix1OSkfxgceiQ
p/E2c9E5sV2UqnWim1MJTgpRd6fzXmX+1skyYuaQmNvgDOA3NP3OhgNGxVispV02/7KosZPR1d65
iQbw+s0UzFHHBmuX7h3yNetOr95NliJ4yJRpaLSdK6ntgKyPvIran5yZUivTJsDfB6lP4SKGZLbd
r4lkl59lyRBsZMcpnkFkJIPmCsBoPdI0wz0OyUy2nETkvGW2YFY5Y44Kc1SVxwqt+wsW4iEol7IB
GkSEG+ofyD4KCsoAPGWGpkP0RS3FxaDD7P3FWekkwksjr4sXWbINj/RTGy1vBUpHx5ZuBsWeD3D7
dA0YEgyVwiYG0sqs5ErRovIBtUYI8i59YxOa1jjbtg+yNUle85lAeOOqYuQ23xSp3yTuUswymI6I
aTzunHjmjC858qcmE4lkRfdX/1fQaKBU7IsZiqo2/LsxqonyB1Z2l+Sdhsqk1zUxz8wO4RE6/ze6
OlabJ2wFvxaYsTfXjSt0II8WhogGlLathLzdYf/WA4PgQkGQwh/dHQb2zEyAI4D+AfvaQWN+dMuU
OdQtxCWQ1vUgaaFaeNppE0elXHG2ZHQBPK5hnfSNcmrEBDE6NDF4shYXbi+MKeJ+zzODRxengSKW
rL3PKIDuQlryu3JqH5vqslSTh5/sgY6H3ck2SEn8p17yTXcYounP3LakkfXL5LAucURGNzIFzLCN
OzcTt9FsNnHaQbpeLUHh0qRmhUa22XP8C/1us3MuaGdMlIOTmT2uhkrfuZTejteJqtio4GAQUa8x
24KFBcyDPsIhPaztBQrZ7R3bvXikHjYsWeoaix7lg+bA156ZM/2ZDsY0LaOHbagt6dUKY797ERiN
vzXj6TKNoV/aYrovsfuVCvWxZE7T96RuE/xmpVkj3mxeRTLv5sRw0Rwns1q5G0J8KNCeIor3vvFX
E41k+36dL7+1q6rfctoS5+F7aZesae67yO0t9rrLBCH0yAdtRm6F2+OFNyA0XZOGeSG5VDFTLX00
DX9MY8Xd0QHEJvXmtwHM3GkWd5qtfGbIZr7mOQSyTwRKkyfzvjVy4HtzMGSL7QhUbmCz3Ae87Cr3
lm7g2lDpxG2Y4vEtE796X03MZkJeg0yQaHUnLEG02SigGshS0PSFuzxVg96ddj3T8jVYL80Gevhr
1nFvGoG+miRUIpK8oRf2V5WBLUdhol+ET/+B9nwbqEw4PtKXZgq3BPUOm1BZVndIMf7HWHuEUdeT
Ze+5U19yIKlBhnJlqtywXOfLjZ/KxWmwzfP7dK+sucAzyE5kGjnxAX3AVbD0JE0DoDRAarP2fl29
C3320PXmCVU0TUkBtSGjHuvHDuMQRo0hYodaVVSg94GObGydlQE/O4FSj97uNVDwFn8x31/9QIGF
YMfw/RI8OygCmAfwq4CdtlWYz9U81uIf0RjP0rce7tybzQvbs3hYCuZH/KfJNz3Hh3/T+tpVhDTl
lXfk6wFYoJFOVo3OxNTtbJrgArxd5RYhRY3PgUJaTAZjgGQuGTvFWFfq4hFjXwkX6FU5zCVwZe2O
ZAlPJyKgk8fY/7AcT2keVHPGoEO9je7d0S1gtE/F0/pPEHDcB2mmp+zJ0gi+i8gxdotFcwPB011w
6VTlk1vijkkZrjZjtLoPF5eoWTRuE85V00CouVcREAKPOsfeNZVxDDMa8Ib17/lyOq2+JK2FF2JF
3ddz4Q9SJZ7GrxSKBCrsUl+napTtqO1gyTdRcBQO1RLUnKH6ASN+fxX1SAsoQ54dbYjnLJZ0XWxp
qYIcxb7eWWNb5JNDw0IQ5nuo9KsZyqpg+Uc74Fm9oKe28Pt7Tp/ux0wrYO+vhUzt165aG7aInENJ
Z68Vm0OYwI5s6tNvR/ER+4pRsUsW21kRKt8mYYLpscbLjn+QyJsxLoDAqDSdvGsuvkcDiMgWsqN3
8jpnkoytrXA4wm3DFkBNaJlMyadLZVCYZGFzvIN6mZchxFLptP9Wlm6+Vjx5M/qKGlmZYBgWNdTe
sa8W+UFMBLphQHZoqwwrLK/Hwd+xk/Jru+NHYILeiqai4KJxTeUOhKOoZOK7Alymki0isd+IeqgC
6HGFCkcqTaXafJWd2Q/GDXm4YHvVOPxOrs6otkZ2EBrIoWuMKqHxR2WFKg+LTGrdL+McKKDRPEB3
cuYK65xv+yS/PszZH1vYICQlLmO/V+jnlFCadEh2A3LOmJ912xFISjOQ1kbWqVJREUVaI06AJEfI
AhlEr/MlC2UJgpe+oaTBrouGyuzmmZg/J3xNYQjt+o12SeTxfnnDwDlj5nteR8XWY6F6yLkYXkrE
tDLW4bCIhUukXWMN1EfcNEn4b/2NrXdWSc8+9JsHqf8i4W2Q+vhnVh4xgIW23V0c69nNzVF2I7Bk
5mdILQG4DEchnUhLW591sFy1Gi+KzFl6KSzRtf2gEjYo7U/WM1egfjJD85AR8m3fmSDKkYjmnsrQ
FiN2sLcNvLUC3syJoCcPmEbUfzasuumNK0u6QlaqwLbpxqmCVcS5mLVgl8E3Ib1CYDGdHgMx4N+S
mxFjP7JC0QrEB0vfURtH77ejeganv7ihe8P0a/synMCZVkMTgEfg8AFy1o+MuiypeO+V/fCKDxng
vEHK4W4QYU1WgbKSstO/n7pj7I0CqGBH/YWIL9IfEXna/+o2rOefdbuFAd0fGzTy6w90lY5SAXNz
Dr6fys9hGp/QAmliCQfe2zZWkPBaC36jVx7eZFz+DB1ml/XjCwsyZLRkV7DbQNJ4kgMM+d8UD70T
0rsqUdaIKnUBCHYNGkFPdiVYQDNQzqq6hCRaG3K93WrOHUQ4l58adCFxu5531R8txWAxK+NKwXys
7sB+JyDRuH2K9iXzarn69/is6XPgQVtqUJc2WAfLV7C07gop1QH4yZjAv6ZND8kYpWndDti634UN
PKKjmQ7j8bxRlxLbRPZm6pWsntd/0P2+4Kl747nOqC9QHhxK3LexqntU6udTjNHtBkyEcUfgCzno
5nBZpUSr6lN/ymtD7SeC7Ta2VJBeNUrtIdZbSgVZvYOCzeQTMwSTEpAJuD0lTWMEmImdTdWlFIOy
I9tih/pwbDCQQzMHyj8FaQIaBhe78XAmFpZJKvHxQcBpFjg3epkOGFgd6dicemBvITAv92W9n/sF
zmFtWfMRbLsfGplzH3S5zxX8YtaJleuHLh8zFOT9DpmIiYxMff/9uBYbMkMu/yzizwwIUi/0T/Xb
5i2RYvSVgCfSZm/XQAddAC745BKZsIFA+lsSpRLWu011NfnDwRCND5sOCyEAEGu1B9yqVdc6nI5N
RhJ3EN+EwwYbX5efPo5fagonwteA4D3LVXKFj/ppbJmF1a2BwZbTX4M+wwwaH0dmvnvCapmD4mQF
A+TcC63wQqtMZYZoSG6SGrPSp5i7DOLz8sX7gCSx9fR1mdSJvBnT/KUEVrZWf9QsGWWbzueN0UG1
vNaCbQNWb+d5pHmFflI0ArYs5pq1hPdKd34ZCoAq+VNIRO2OUE7TyBtnVXZEbKB59YQAPGXNjzdg
oJxMAeRfhoDNkqRO11u+oOuMbndMRgvSdub0TE6C1GclLxCVdLlfcmYyhEEIyj7qK5F5yiqnXs6+
++4McQ79Ih9f+LMXybPkyrOL6hs7XSyTOen63hlt2Fhm0uERVny2rk+bfwfg7AR7A9g2rd8UgstX
KOrB/s8h1BYh40JS8bptMisrbm4PDDw7k6gWL102xrOt8vnXQ1PdNYQ2ydbIv79h31TQ9OAh2LWx
1vILEaC+T0RwTTJXZ+3AA49KuuvV6zApV27r6RRG0HQcBw2zkMjh2/Bgragd9Ahtq4dsZR2XSNVf
efF1nzaWgl2Dw5Afd60DA3TbYIzv+ssfSjawdwe41DymJcCrAtzKvDIeV7u1qPPfrnwGwkiuLbXj
bvpgyvi4qmAIisJkkXqxQBxeYXTSsn0vqe+Roe3B3ySP7IoyganFp+Hx/0cIAilFaCmwxFb6vy67
27LSH913sOTtbfrFgET6aag9wYC5gPwag1Rj36Z5ec5pSYSHralAfapEq0tGcyBiym5y70SNrjwt
jT1VpHEZkOsYH1Oh3GDD425llT1BAP0hcXiD4TrutGclVmy+rIkaC+UaX4ZdntuNbvedPMBpT5bW
8RYpmxY0g///MNsuPcjsZHrnb8mgpDEfqnquhIfAli2X3/tZ9IiY3ZbKFtGMAMMv4/sV2RGed3Ct
Ctb17cpYpkQA0QpUwHNuZHNcrQStD9ygbKnCs8wlC5bXE9nCUbtq/eQoHvuxtU1J+T0OC/tkqCzJ
vemFIcsDGtTOkXhMI9TSFh+IL77029/hovksfgrXrJ/EnucZ142RPKOeVSWXoFzf4LTXlNBrDtnT
n31/a2P/V1Ztc68zL5uoBFi/PGjHGt90CObKZDazvaKYX9TxmaOWKfqKLliPjrudj4cvguSKl4tp
AgsdP3qZQcWyhegupXZCrGO3asrJIbIfDiEf9iyA0CzAArihCH2HsKbcC1RMMmWeprmlVxpkSlaP
7EDkcMw3ClLIS51eYSnLM5XIje7okLHJhd8SU9SvOTEje8ux9kdXiH8XGnhTzdH0veHiqDxDPlNU
UntipKLfKR+9e/60sM3gcCuWw52dLwxxKGV8iNV8DuN/FRfy7qgGDLcNLvwTpnlbeNhcMWVpShvW
CmwHl6M0hoDO0XbIDn9nRHqQhcejRXthKqIx1S4alHVz2Yk/EXVP3H7ZJmV761w6ORb6fnmqNQut
hmaLtAWLTlkmODBzDIE8bP5qSeAuKp71YWDHbWcQ1Z7526PhQL4KM4t8GWyuq0d/2DE+GF1aHlTy
FfwJQFLek3mv/SSKiMm4bcyvbuq9LvNMpCuVtVf1c2gHOes7u3bAYJi7BUn7WyGGvBonzXoFXubT
6SDUbs79eE5UMjNwoIcEmZjFH36WtdYI4+7gCxpj3C3TKYm9Y3CtiotZRwHggPUxUr21J11pwS3B
aQVj359LHIWkYtOEl53BhWkHAb/aK+j7oucPDOEsmzhkqPiY5JfkzXGjDqHqz+OquglXd/fc+eIN
tZ9HeIw2uGz5TPsFFw79ntmGmqdU0fXlNMy0aH5fxAS2SnNljU52Zxua1GPkKofZyEPq6zQcw2+L
FJu7G57HBaEekFq0pZY55ylM9wDrdNRbls/AVm+WVAWT3OHwmHYuCJVfUY1zhAF7TFQLnrbgfcML
xjulL+JLV6N5YybQHiOx97lKXmRMVzqdPmS8q4IIxKYASy+Rzfige7Zmj2RHb1KI1hSxfBy02PmB
qaTHUI/rta5CWBuS6GhU31s1lkDwBg+WZfryCYLV6ngs75NVA8KvYSrsCRhARVTlGPQa1tpYQ9t5
gRWNbREKMLpI87ABYC0d/4WtWbA6HiSqNH1kxGh1tmdLPTaXLSmiHwO4q8hYR1ueLma7DB22Si8c
DuusvmNi6+tMj111afsg8v0JlFJGz25VaAs2JSIHjurcB4GcZFiXOvHYBN6SKtw6fbpnM0hB5Brp
STKa1pJXrKti8qWP2pmL+ObIboxTGaIFWFDYsn4g76mYo/S4+L+THGfQJCHtd4EL07Eik5hi8wV6
OSX0BBRLHfe9YHTSSt4tzUhHy0RKLECC/tZSfiFcoNguhk0tehWCtcNhwy+PGOqQd8i2fCF+grEf
5TvrtD+mCsypy2AIhl5dJm8JGyvT/okeQsf/PqZIDUzgobbZTRyzGbS7+22xpWr0jJ793SCQmyUp
DRvElubnUme1Pgw8jYRICWy9x0flpoCsejYfqBby+2VAovQb6XUsi7Lr0kJ7ZT6ZCkvWJ8ZsPoBv
YvQaP13EpXvKakb3ACjZ4FFaop2t3Qhmhwi8bBAs13dkOw/0/auLouiCiACbM8v1pXxgC/uptRed
ZuLmsLm2O0Q52CbcxXarAMsOfLfngIFhqsR2AojZF06pjyT1YWaNTvk4NwBsa+SmMqctInVVz7AT
ppnq40U+yFvIwLEbbcgDHSnVc4jVsNOOvrVIk1fwtIo9Pyp80X+w+Mi9HrNkOXQHW/1DdSV/TfXq
fryXplv8lsDLtkFPDiZym+NqsZu89Di9FzyzI2fDJHQIrsdE/7GYzpfzIekNNGH8gQVOSEFxGT7+
vBgRbQxaAmz1zw75GpuwBplXE+QfSJL5StYzvs3QOVU/29Nm6AD4xI7LNp7FgxmRG9+mgiS2uAcM
IeHHg3gtipAZ+5gcsboy82brkvGbShCFNqkYcDScgs9IWpjx04Y6Cq35KqRjjSOt4m8pmRcjMEbV
8M3m1av4OCSHJLnSYMotzgNGfd0WK1Gpia5d+dBgCFoUFzSSnLfLOOcDX4eODhL9fm5IrRm013OV
cM/2jzCwapAm7UeakfVUrpIM0EONnMcFdsi2s0aBOIxhfT1vhAPN8tcm3c2qYU0AW0i4EQ0yqbBv
/ht8ujijrxUtdiU66xU9jCK63gyqZnDnRGxFl1XwRUILICYfVrk3qk20tdjwZzb7PceD+EStklbD
a8TttivvHI0ZOrplGHib+P8NDlUn6t2IIhSSsfE28DdfLKJRrm2WMcfnFvu82i6HcJX8MuLZAn9m
xTPguBBYCs+2IxIJE4r4FjWUqA8Q7qgPCALzbQ+Vqskac6S/ktJoe7+1UMlQHKwY+rapaaSS6bO8
qp8DHAiKGtD5gVeALCbswP8Dxxobd5PgOEYgYwnLLXr6WD7gC4ScW0CXFFiI+/d0K52ZxQvokxll
ioyA1mCJiyJUEK4C6X/gbzUGjKKu0kZn8sRqRoYmGI3NbeC3FVIvK0eQtYU2X+ta8dnSob+17JQk
+8+yZvv68LPZ/YmOuIm5L1OsTPayTFYfIOYF3QGB2chHiZS5SCBrhpLh591zPX58r0kKpDnZXirk
y1iBxJHqwm7x45p89d/WqoC7oRVDZ2o1665EQB1eAPkUfYI82toTUKuzr6nIwB9KDvMffsW6YWPL
EES/uj2AkYZQf20od/E25UB/H+TgNYVi+0ojeSu9DSrTCAitW/SdClbfZRi/aXItvefMGNJcmOVl
TLXd2G2aRoc/4kv1nCb3cRnSPq5p5FsumR9CKzgvDD8ZacUYaP7eH0CrUuCD4MxNst8InL9y6LVP
cdnJ9Q71Sh9ReJuh/2cuDOpYLcSUVfJU7ElRfdhqWhJRQtHhpNq6go3IaZSxQ3C4lVJxmnGIrpXY
275730TmORJsFBOKtiZA13ahLXWT0EM7vq8Ql+DjN2KQMk8Of2UKs8GDHK0vYab164EmMAL/WBhD
08lhlmKjDITXn383E3UaFlpwuB11KCig7a9TWVF3mcsANMpxyyzg1vAy0cA+2+1q89h9rvb8XjDE
9vPn/BaFlFuPXdbdDM9mgGAesZeG754nw6xD2lAoHAfUlWlqVnmPed/sYF5Ci8K5G+gHQElwulhO
v7gQDyhlo/TCSzwh8C8zrr5UU5Y3ulhqBXUIQmFVRe7k+VJ68eDn69OxG0+ON9/OfO8Ub730lTvD
8jJF++6OaMOMHNNKvMPiiioKr4AnXVaZGMltWCxB9SFl+RW/DGrd1Ftx6EDTWrz8SxJBDeyJo7DE
vh+68qZxRp92zm5thrShtJX8BUDdBnJlgV4RotlQgA8WXwQHhzAl2hzNne0xj34kPfuRNYbzEox+
dz6MHExM/eX+qaB+n0HTuwFwlChYQ1eg535wxKS/GbA4X2bTwjsqrJ19an7/u9hw4ghaPIJgHln8
ArK7cLf5bQTAgAPxudR/cSUPt7zD91aFcHCoWoby8CSZSIP8eQKNgNAlZgPfUF7od8UUriiBjG/+
0TVeJLPOJLKSjm1YwzPy0aLBxf2TnA6lu+lWKKfg+VH5HHFH+I4uol1Aj8iJ3DAwBzL+q6gpNTLu
CVZ4ebxLn+jWBDAoY9JU5lUfMI0FtDsQxXwzeLEQbqlpY5McoIjOW+6NlQweidmhy2YH43182PsY
BNhKX8St0Q6yPg/edBDHclPvUgmS0sHRB0ydymEBZKXHk57/JqZ59++FkfBDwwHxFm44tz3KqyWM
k1FB1LDLMuX8JMhrwdj9Dw54THoAyTw7b72iLJMXh8umZG4lpfB5LHBhBgAoPdWEU5kW+aS67LRw
FO6nPBZQSunKdUOzKyeyFeA5xgSy9jbRGbLwLbj1fxoMsCMl+Z+XyhW2+wWfjRuFOoHYbZUHgdnD
SYobwbsyBGJlcwmYJFNcGLthcZBjVkZCaeQV5RPRoISZ5ADYeJiseCyQOOf4r3foexSJcWlOKOsU
j3BgLEltc85EEwcsIpHV1rsUVqQ2LjNva5DXSgDzUBeBzk5c8jfohAgyqpKx5nOqs6HORuwDQSWe
z2wH6MiVvty99pVWv0b4oCOoChRSaKwGixilraopiaFx90nkoUWCqd4j5YLS1ywxOQhO2AfhmS2q
m7nlkl9vBj06CnF5BJb0hYO+AgxeW0iHnpuSBmxRJ6FH1+gsqHQTVsgX1kcbTrQ3fF2IhxiKG7l2
Oqlib6MH78xAp0ythCY1Rg8ubyOXtBi/Pm5bYmiJLx3O4skmgIUy9ruIBWzdZWLE8X6q+GAjWHDQ
fiMK3D9hJJBfwSdvX4yc6SS5RuSwe27GwSK+Hfznaa2Uw2lBqqp1wm/4sOwJTZIFOyUq40xb+uZ5
5B5GM0Znrf5RwdFWrQU+6/dNQ3OtmoYtxaoTjRb7b4FdcL1a1/T21JiAh0GDAGTsLzldN1RbXmBD
Byb5SX0IoRXgnVvW0lt/ircYrrD8PoH2RuT6a4IH4kqmLB3VdnldrhdJJxn957/cthvEYeXU8h9D
gT/H+6e6RxlJ3QHzJ3Cv3CBDGqr2BFuI1Ze4pFZct93gn2aF4qiQoZ1J0QCU8ZiYJyyf+qR2HMeG
jXjUXXcigPV6etxaAzj9eiTGxaBLMz43e2ybg4TGVv0j8SJbNRNaoH4TCoM7b/a63H/qWSeRFBrg
kcco4DCM5URWynoRTPxTgKi5kWiC7YCre00zEFJB7U/TdGf+ufdaZCqC/qB+PVRy85nM0TZnQOF4
reS5nkIpBC1vG07dTRjnTVD/c/PIIiGUgsM75p6w46uvqUMC7SBbN7xbV029GRUJRCR2virkVedg
CR+JHbHePzww/SYPdBxkz4crNLPwBpTytNqjR+QygEFZizBm55VTZEkN0knEzml2kV2eXp1IZZOx
ZqDjMK38VIr/Ll3afr/jIBW8Fw7U/RMGdV4SCCCHI/1WJBov7d2hi5SUhBsYfP//eDbt/5NKZlQ7
5Sb4Hk75IEh/JfQSOZws+e5CV+seULpl1pn++N849nQKkx+gra0v8iMTx0BIs04VNzqIFOVQ7QL5
+idg4rNdSiwZIHmFx4rT6rttsKrhtLMl9AatxcRxzjbWpFysKFQkABE3zAODVrQKIxBBsS/NS5OK
3EwGqWbKgIcmkSbMhjwvOad42Gw3bGHQ7JJfH8OSy3twJ+uZrgfhhKNsIVoNSalRkyuORQaM3qwt
HdVAoPrw53Ga1Wmlvt39MXTP8vak1BnOIOdd3P7HuuEbnjZHjlwmVIkHFVE4IzGPvs8rrMFEBzR3
DsDOowgugWrO1f4I8ofD3cybOyT0uuZVDHyHboxVWmRHeh5V+NHg/46YYSCNf5yKTVTK+6yWsSht
99EJXxv3NXi2zi61zKG8COLTDQI+ZhjdkGxZQ9//MYClN+8jTIrLItPTox9/QR2cMyc7Tdr4hQHq
KGHl/8U00Ea6xFyDIMuPZXX+v2p2jWjJoAU/efsjVdhbCLm0rjuBRW8h/wrJ0DEhl7t9jy5SIuGm
bI4MkDiLSZ9/Lf9vmg9yAnoxgGpihsQ7DIh4X32Use5j+zrHgGd5GtSN83CW6D1dl416jbN1vVmr
fNHDtNwjTXtp4O0hygdc0jZDSQC0YPfQgaRAnpdx8SPxBhmVZ13/ksvBHX5vFZdSS+/PwKLKrTNG
xFNZK5mMHypXrtTrsVMcSnlbKCLcvesx0UqzLrrh7kCgmsqVHZCGTerJhus/xivYUGrcj2CkrQ8J
TnMVs21dExoAGsSm/2PEOop8pjDYu2pj/nyQFd+aaA/CvSWT2QTXsr08pOQ3IbmH/9NqH29Fnv6/
UgDcVAIDQ5GMY33clpyDi9HztXgXlbXNjE0tJv3IJp4pm1b1u/mevxsVrCZklDJTJu0dPLBf7Rsb
muJhVjgiuafqTr5sZLG1Rd7653oD7ypd9kee9kJqHqnPb6jwwFTH3qMOads5yFIK23cmA2yHQtJH
+iergphFL4kDT+lA1V1PicE/ii3IuZjGW1onH7SIWoCocDQs+XwNkWRfj8U+J69FATVHRQqSGC5x
5I0Xc9Oof1SELirU7G4PU9fkZmzm2CZmFm10lSOJgjhYg3gv1R9CMYDN5m4LyV+OPl4iBOt6gn9k
/ir1U6c1XQse9juORLJzVFpfOxNejyh3rqiEMr4UIs+quYjXwxlREn7Wi00OGg2Mjs0TvTuCa+Ap
g02R3RXclgBHiAMVyPOeZvXysFh8klAY2oXLLny2qU+yxj1KhE5krLdXtgexhQYQvKrMt0gWjxyi
y6jhJvjI91FjPA9GSJ2Mlo8AqfZCSEIzUrRhOU/o3kxpS8O2KtcLUmO7SKlbJdyg7rNEPpEJkYny
WKKuDiWT13u5bttBM0KIbLqIaF3NZ31ywpP+RFkWuZpuRKdof8gVNWYVyZTtPtsw5oTKMkW3zX0W
zpnDAwG4la0R1grQB/D0OF+zEiLFZtZea1VDfiBPpIk+H2Ofcg2KRJkCvsoRUzsb1D6Gw8f9Qs3g
6nYyHvDUmnGPgC+9V8pdrr+eKfiaT8FqUU2Jb4gQBRPCjvOeAtZ2h9pzKbIHcCKahDjk6uS7QH7Y
riGKyhMCEqjzXSCVBM+Y9Q7ywErFsQTcqBsqjxXg1xOELV3eD7XN3xkHS9dFTEz1gyrzj8UDg3gp
NhCTve/WH6NIS3M3YTIV5moHQ/Mk0iKH8spN29b2RHITpAilfUUPGKyn0EoHPFKDx6LSsiiygEzM
F4Y3Ak+F9bhaCbYPT6BKYK5Ej+z+cmVprNLY/8SGOr4sh12BqZ+uz7h+DzFldZJSOoJlTP5D+vgA
fZNYUm1MEpahx8tR4PsqCOpB7BTKT0LXswHbAc6/Kyz9iFm3zYldwmI4AdvRveUMH6vvX5aTK709
KR8msjt8vrJdSss8lSX5M2pAMofPn3NhxBgFBjO6yXt4aB5a3iyw4K6Qkvzypo1kKel/mhouEpOu
rh6XZW/y+HsnPz9c4bET2/6J3ZbIzuDpwjgMjR9iDFeTdyIpar2rfnD5+brCykieucom+/UK1+h0
YNyBeT+NJDWVYLwIcP+rlEtBHdym0vGnqXfaGbRKBnSdF7ZEzhZL5jq6JzxpxeY1QjaBsPRA4nM9
gLxZ955+fY/xfcp3NpSK5qVCIfpH8LUcIh0iVa+9s4bYIVlS5hYuGHX6lumpQ9Fja1O0ekeA8E30
4a/tBYid/rfXHNNvMBTjkxrzK1dm1uoZuwrfFXFmJYHxqoFQ5XVlhYQRAXZP7ML9/OncUAsCI4pz
jCr5t6rOe+JNGGGiWAw26dWNspecwcxH8iW3TZT5C8osSCJO9cFoTH5LObm26Ryn4KjQjh3Bv2Kq
+3Fp30WTecix0NnKoO3iKJ2CogYGvGehich9kY+2zgvaMynqrx4aoAyhjOryu+HaydbAFuETQJGX
KMnLjgnclnTY5GbIHbLLN5DA+FUcT8u7WgYDKbEjhQsRKZciSwMlTDqnJ+ZlvfuBRdST+KMiHEP3
uYneZe1/V+0SYdujQvg6EL8UhjDeq1BkeQEpAWKUcY6UVGMrwGacavJEsqkydlzRgezXq4Zr3ImD
mJxdFJqHHT65d9hYVJzB79CsOpRL3xUNNwZ6DghDZpWWW1fie+Kt4J3UNZjgo1hrrFVZ+0CpmIL8
8FTDvBGbmN5qgx/TBrn9ofCd3XbuizQBeSqFzxNVzJgcP8gnksov5qV8HZFA8WtWPIZOcbxiRdUJ
49Em4FT6jLOB6JJnHZzAI81n42ZxbNGgX2nzks8+L77zGnxbpRIr24v11izf1r/Sm7dPUk9oDOh1
adXsTKiQT9ojFealkecRq9IgOHk9IbwWkFUkzbolxlJihaS4prPulJgRssl73UNO8nfmTOX3ixvn
QkDVbOTDg8dX5nUnddS+5C5suEoBicwNwfhsX5WV+dniSjKQxfXTSSM94GdvX9lb9kFA7FL0xCL9
vubr9V1TD+E0zMA4DqCNn3/63tg6UtxZGn5czqbPp6cthcbMg3IVUmEGPdkl0APH3upwMvpvfceL
gGXWSjf30i30UbcpBPRxFU3SqxbcHc94je/tJn2oDa6mOBfmu94UOljLXxt/4jFXRG78V2Pvb2+y
eMM/oz0nlCxDqDY1kG4RyFXzcKUqOd6vTFcxBPVtgseA9seSa3dujetRop722eCJDSyrtmgifMB0
ygfaVD3am03+Funb9fO0LndIH+CMFbZmP57UNuFSFNEAk6TZTSbTYkayoGgD+42ypzZOgdccU7pI
xX4lWBesqBhiOZK3ANVpzHZbXLE2nmR6edybRzQ6GsfXkurnNhxxKt5OYPWy4AdfLIZoeGrc5QJO
J6PYYdYqyJ5SnromEk3T1VSzF6yYInom3FwiFsF/ueidoMEwhQYxk+kSfIKv97HsJowmTshNj71W
RrtdLJK5JQPwb5CL6t2XZTH19dlsW/tbEvgNRGoWzXTey17kM4WivKBK8IAZSkFuGuh83l+7QQFd
lnRa6mpcKdO81yqvwR2yWAM4IPFbpAi6FDKtJd5+rscYpWymIvtbkKE3LJgyPGV3M81eIRQTYL3h
kqDMJ7zsg4xW7oL9EIdKjWTBuIn23ERzjvhTnlfNDDjfEcfZw1iEzT3LbPmb/27H455TfWmGq5i9
bTV7zPEbxdYjjrW1tJzAHZfGaAqtSWQ5/7cHd939bQOFUQy+w+XXVHHTV8WuLxl7LPm9YSw2SvML
Rpj0/QdsUkLXwfpck/9BiwE/m/1F4NH3Dl1IzrQ1xi/lxEDlEV+cbhde+GojitnfDGrgyxHQ3KUP
rVUMNqq1wZT8OTmvNrKF/iseQbPTl5Lw6FxX+6akXMuBi6AkZfL/3uGqPTERc5YjrBEhAsVkvU54
NE+lrZHZYP1BDi15Dy7Urm/dzKMUWqeq4Dmn2nkav5TaLjssVCnCi+grzfCLrLyewxXitvL41Rwi
jkjTRG2lKiPwEMtk7H32TEqxwJRHN9HdYeYGNhOEf7oeWDL3AlTRA93adlcZB4zt87rBTAhdsMFF
dQlJ6Km7SbGD/J6T422/lHX81FqpCMV0puCRt3owdszcIYN2/utGyg3xRltCY3yjD8B8Cr5XCzMt
h60AA1moJrQsdri9T9jO/Qdx28WCpdk6UI+zTbwv6yDxPZNU8eQs4A0KmRC1zfL0Dh8td6rPCtrb
3IMM8Wo4uuayqVjx6Az1P1bsQ3znatsTOWfV7ld395txn186mwaRBXnCDRU2KiDlFzmFkA7qw4Gx
GktDv3nXDZGJDYohIWJQJSo7i0ot7b/JjSy4+sYdmO789hKFssKB6sIl3CWHgMknw5gMxRUJnyZ6
x7SHg1m2IGDtUx1MAjVQpC3E7nSiDbWyEAN/pEgMeaJBau4/qmr10nKLZZthRVnOVPU8f1MMV7Jm
WTaUT00YKxt1zkD6pbTz1vG3P3zBm21GrYjzJ/1fkEXe+r8IUQTw2CD45eVIXavOeMIRUs90yeUu
3zAmpdd0xN9A0B5GqbBffslawrE/PFER+7+pXAflo73hpvoPfCpSOLuU3ZaJ7xxKDOZVYCk2KeiL
SU85AEbegR6SqfP+ZYtmAT8i7xtt/IQkr+UpQqEoPH2vuAjlFNP34fx3OPclyNwYGAy7cEuIBR1s
bPJjxI2T9OoyUVOadYowMC//onloG835orkYXxWkVOGDlbYG/Jd5d56ZeNrZCsMAte6kWncWONy3
K236PTDTwWMGCC7tipIB2THf4LoJ+IuZ4PU1b04KSsWcwPFGptXdm+4QH/CBRG6XzHm2KBouuthX
mch6ATbHJiew3Ous634ixM+BD/kVW8qr2hO4toshK7AHa7HfcfnPtS3mX9+V9aHA3KlH/wU88rwZ
EneHELBAFInEuZocCCnd8gpuUiPyN9Y7kPFVBv/d+445fpF1wixXzj+Vjn8ZJgH2MY/UHUZ07PAI
ANlxL8GZqmj9zXIuEOAxgqseOJf17v9KYMYntEGByjvLlbf14hcvYX0wVLKqYUWHkCfTw4KCHAP6
Wp4oAVZVduhaSfhIzP6m3O7ozwlyL3MLuuJvFCPDKEzPGabnMGlfY8DKHuC6jsZ56tEbzF7Q/byf
7d7Z6HbPDFUuFnPUtcebfkeRE/j24KTg3g1ELFY6dT1Akd63OrH0o6WIly2JJEVEeD0Grv6shZwJ
f4V4zeQM2ZtLNX3rE7Qoi81s0uSU631gYVOnEjm2a2VBxGoeEK2L4tfmMgxu4dspvyhKQyYdIsc1
RYkmJynjpfmw6wIW8YQOnIEJsiMM6ltT9AGNm8wdchokpUfh6YUhIY1GDMIjKlWWF4+UEFdVNvxl
L2A+mlz9YcE9yHY3BAYDqFKbvWOo/ruUX9Sbqu+QaOppFngPTTKI06l6Qzz4OzvsT6u4WB0YOGuI
A7IRc429QJ60V3UESIexalZXAePL0PgRlhldETxST8Ea4mzQ/mGiw/H1Tlw0tLA/uBMykICm5Irn
gdQJt4Ez1qzjHAEBFgCIfienOHGyAu7bdBg/hclDitH+OglgAyAcTCguB3o9wQv4GGU/jvAyS4If
RnmHWnXjXIqbXJqefxvaa6rfStjvDDc22yo2qJ9a6sM7eA7LJwWjPZ1SC+uKKMCmFpY0V4HPxs/l
1V+9zFwi9531aXFXvcFxGvw8SLYhQIc1WnBrPCFKRcbAitrrasbxF2GA5284zLoE5KBslmTZmVcX
5rzP/tMDXev3TCOg2rN8nLITC6Xrn/bAafTY7ZAWlarE/Ac+dxGEysSaQPU0ItpiMyAfscsTwMl5
FREaMyA51bjCCrgQMoF0Kqz8CZpU+lmlYiyYyYPdVoxfBnL+NfeKkdD85J4Y/X5ddc5O43RPVPE0
e/To39O/wQoYGzslnCdfhgsEHZQbvQ1V+srS9TN/cjHmshz6jHutECFneY3VLyyjGm+pHLeQlRvT
9Fur2fcXYE4P5YP/fd+GMlwDDW5Vn/rI4RZBK4htIsji9/c/Omfkeso3+LWlnTz3aIckwUxAWniw
xz/+bw9Zwbyky1OUBrQld1E2Tktsl3+QmGnz8WPrnsAaaAJTl9kp6J+qNVTIXZVc8R/YXnMjBdyb
0+XGPK72yKOfjbs4nqPnoQFknbTklYNt1tA68A/TB/6hAj3BlzfzFsUGLBm764Xtjgu1Sog4WS+a
1JH9yPMRQniCNKYuHQjqSzEPvFfsS8ELdSVV+1GJiUQM3kVMYpsw3VCRPElgWbXbhKynA147/lNN
uaDuzpKa2m37TZgOdMAXsT1XDaZyAt9RHoi8POpyjNilGLr01V/98XSKE7Ax1yEekIXziERgq5f+
Qz3Gbw8UZX2CXz5auBoMbkXeBY4TTtNWX2wpjRwysQijFaJBH3TrDASXsymXO4kPgYbwXCfp5vfx
lqbQwJbDOX2DVyNM78rJk9+l3X62cmh/ZteFmlETBVR2wa19SzcNKGE+UgZmUPozXlZspQWvbhjk
K+j3z1rWNrpHTI53kalf8v7TgglLz0IhjYxFuELpXjPTHke6PfWcaz3ZEvvor3tVyg17fopHvkiV
joaI1G5jlM+a0ErXmE4oQ1Dv+kSdKKSflmmHt4e+zQMZvoIektGoCwisK23+mknE6ccnoPHB+wJ4
wn67mXrnYWf5Jt6lcSc6Bqmcc5TNIf3W7NMHNPbcosOnY9RM5xBqBOcdtPCInODQQNFwJHV0V4w7
fCclfHliC2U6WYZwD1LKz9irRxV+4I0AsJIMDD+FTosnu1dK8iiUeF1YFFs/IwjZmCJJT+TGT4Zf
Qw0xooSOj0JldCE/021shCN1yhkX8I60LVD3aMtZxUaI04CaNoIfcKcrJSD1cmmI5W6oetbfx8Z3
lCeiJUy3YX1R2bkj+kVmq/UvrmyXCF9X/omJXmu+BfhVliTdO8aRJ+2FaBSy7GKiSDMEF/EtUxhO
7oGnfK191LktBgSumj2cFDfPgxNIxD7SSH7rG9FPrIB3ZpwmSl8dmZOw34iEkH21gllwhvJeKn/7
d/7peUPn6PEK4XSv4Wxw/19kzXVaW7HmEfHIQ2nsy0Ewc3O7H9ijVTM46z9Df3ZIOEjCOs8PCB7V
KNPVki1G83wndKUaldnDotzqcb6wieEB+vadpysFSExm0NdvasYiWa+z1AfrMe6zXwWnpGdxokVH
p3z0Cd2jrCifZvx+/r2AqudCRvEXsjKipSO3gaebM3G93frDd0EQK8xwU4BI46s33g4T+BD0pasL
p7Q56dleEHRXr78yTuATzCh1dP1jt2vwgw+lDZOP10B4Y4pVJWY/mOTa3O1H6tzyI4QNHKo4sw3Q
GMPAAGCIMwX/sZkpskq1xnEcZnwdDaP7ab+5/XyHuHIUeGbeBOe1apsy/ibruvjXRJiB9cHf0Wx8
FXEdditgsjdT8Mh9QK4oEOD0XetWdFG2IDvpwbdcXGcuTG8EfnIhfs6xJ/+TBSx+3Ks/t/aIVJV0
Kbui+97qSPu/E0uc7p1wf0Kq00RYwBuXxDJm+QLG8ZCYh0/IcDsLxfkW0BZ2c/SaI2xwzqOdNGo2
DcSWhya+n7+i9UNHm30yy85nAILyJoLX+dAT8YjraKjJrSfF3BHp/FWAF5WYpnvvIf7p5ctDGN8h
E0nH/g8UvFy4r7opFlabgB9lqiy5eNx9OzpIwIN1SuEqOnqnet4AmtzL9EOgZDneh4NJOtZ/TD40
m3SCLaFU/5bUfjYGeIX0mAFWJXZJpCIq7mx33q6TMHyMkIcdpvcXX879L2omaqugrk62Fc+9WPY2
pkxFQES2bLGPulAsWUqdG2bKzw2m0zB0M72gFt+vqs+T1PqdX0C+ixrPHEvhULEpY2TExf3cCuee
HDzmIHpEERCZXnK0M2iFojbyVjMbrTJgJA7LPYRslWym0z1nghn46JwTQmc/aAGrLtmc8Q1lTykR
g0XedLJ/kCCWx4tUHYZZgzAWorepJZcvn7tDRA/eRcWcdS1g+CNQHs4jz5+gzGwWtGmrdwHtZase
s+HCRfy6DqJ2UL1NxQz7N8twNxDma426TIFFpa9yptMyLDdErzDHJEtNV2o/h7UYvjwAQBCYBj6y
gw9dXHrE9qJvbFEwhVSsqjb1A/UBvliZK46VDFnHIf2dYZGAZnsnj4dG/HRcFRBhi3Vih1tICj17
aWTEPLpTzjYXNc4FdZRExiMc7bTRYDwI92HXqhdFKxeayhL/6LTmyJRsvu6MmCzvEGFJJrVSrUfd
SMJvjpSs1w6pQBvOJZhvggS51GUdydwPiXHJi/VtS+vuOpbWc4VFYVMpjgclGqVv7JmS0usw2RYB
645OuYbZVpRaWCii3NR+3GUzmNhgPT10nkBcZjGIbR29Xh8vGzuhobXQtWZSYipFbCzVutjoKX+p
jj1km9Pm8ayJtFHiO97iyVPMOFgGerk+TlVAdB6t/shM8p8NcXaIQk3e3BxJMS4tNVke1hX/kSxu
IvSRH48po7+L8E9wpOjvNOL0zdinE4xOGfiwIziWPB2LsYR8a2fDU69jwzqld2Nbv65y6/xAYIiB
CTyt8HmQtkdU95BVBvsUX2vUYFPeGWwS82x54k+N/IX10Hc4BfekW+GnPlrsBqBUXJprY6hED5l2
viZDgHYfvVW+AeMh4HjCH0jipTlmNfLsKTsIOUpZa8+5VVJW5YQYC7+FGufznXvtVHGDNLi3WKiQ
JgKp+pIe2C2Bp/q1TIDzMvCy25SsCzNc8w0KyODtiiNlFtw7amU/OcSeGOnDdmOzlgFUNXb4vrbq
UM5G/7+QeltYq0x7JMkMC0JoWO12bop+xmAWTYoA5qKKe6dOsuNcLP82FVrYHucMxi0qQ1Nk7Ydv
JFtldFknxtxfZJvjq2E2JVqyvb9nwN+VrZsqvwHaDo39VKfkG9Pw6Ko2TCEXm3+DF74gVUf9LHbv
+QzVyXbbInQxad7heQu0OegAg4W0APvSOw9dIJuIlngSwn+l5SIEnP//n6SexGw7OpV9Bc6gY2u8
5Vbc4lfJkd9+SXoUCdl+y3Y+0otR+bafyPxXlPXl+p70kSmYEoOIXLQHmzFr7L4DICQFDdzHacrc
uc4bPHGjN/olDR5rlw0vLaYx+yTqtPH/WKogLFAho784v9i0CfLngplHSQq9dSES2O9ZkiDOOksP
gNgK9fjdP75N7Sl4gPU7SVgSsD0HyXlkN3fGcwKQNWFClk8wifntVNbNCEKcSmA9pShLsvG94D6I
cEhnsbxspLJhUxPJM2hjMqDO+jzVpF0lE5rkskpv4frhuoQEOzddsljeFTZIkI8SZwHDO8f18uCj
MR8DoKJlOxVY7Pbg9GPmvSAQjWiNZ9+ZVvRRPhMrpPbuDV0nltRFwTTwyy+UZjpXE9S86rmKvofm
y1+3l6nPXSW+4O+ck4K5hJzYMR3NKl3DD7x+hfNH+1uTRpIz1OQyApqYxPclZZvl/ivZvatI+R74
bSTRTEXGnYqDXIJXEZ2QV0uL1mcuHNQLYvsvLo4MaS3ry9YNgTUYAUy8fzX8J7IZxXXXCts8SB3T
mVMeYYThYuKLSOroA6KHQqXrBlxNqln/fQzjease9wrE/3tDcFO/7jTtKNuc7rVK0H/j6Hl5Ryh7
JumfNZzEpS64DW5QlSopnqfhIMBFFnMrDnw2tL5N3PzLs5d3cNSaAQOuI7nNgISm1jukDeUyk3pQ
MmM4EZc+Yr13sz+bOr9QB+BGH5aF2HnCjICW/SVT8afhjRv2AhedZ/JZJxUgQYp0bCVRl91l/zPN
T+E/49QMnO0VdOAp1dpOFD4lmJR0I2vAbUXYMMugGAc6UouHKwZGxWU251jHXE3YOI96KcMrbbQX
qN7e9McRTO5awj7Hm3AQJmsBsopkV6oomol/yfCQhbSHxkJ1jWvBotKN4cDoeT69Xfp1umm6g1KQ
mTpVXMSVyXH3mR4Y7KQJECKcVEvWEpW/t+m8j7MijIzNC3aOXr0vpc5XqF4jP+vtQzK9uBy4tdcg
KVYGqgR7lat00PsVCPTfWhy1QVThd3hAUHWecb41CeMnv3i/2ApX7X+pwXR2LRZljFsDyUgEAq7c
DHXvox8YpU6tiaPDq0FvHnN81HdmFzJCEbXSEND2JSOEWrojXWcBt8zRYkIVXYYSYdjvQPaOAFR9
fK8YWa8sbIMSY9JPbbXL6Qk382n02gIzEPleGAk2Mq/Na2Tfh20jMdQ+tNm9tkLHD7FuKAr3wnZj
eZnQG4LU6nc5qtTq+ZEBc8JZ9o5K5bfhpIlK7TehJQaG+7mGYYOAGNQP/5uPr/tYzHqI3s/OxKZg
xqJ2z0jBNJGuXYELT1sG4WikdUgaN7DCYwdNOS9St1IAksZUR7UuVPkvUbnpWyrFE0tQ7EQmCM7K
ZhXPkh8Mq2QETchbzQnCRWPHB34W37yiZ6mXlIlQFREgnxRZFDqmHUtr3GXxuugTJApE8WMCEuV0
ydDIikU97rCCbAY+UpBH7UGq+9z5ZN4qXkU1v3idfAFwMhavgTr5KAjAuozqyw2P7NbfvdtZah1a
fsr10wRsNkluGr61/ZsE7MuTThCVMNF2hedztrG7SPCQaxvm3ZF9pgyOn6KEr+ePPTgzSjrqi52N
jnwDKWsXcGwoxuLNAQ25fZQnX9VsjZyhxYY09rUSJGdsY05Ig2hhDKGbuQGZndDDagMNtNnEY4nY
s5t8GtYZD0GU/+D8mpHAzXnsemH9y4yiUiiexNSegzZjSMlaJeO0v64QTIxzAcWlntGBbLYn9F/E
+abPJ/gNIzDff4dZgkwroQ0BcCYl3uuT+Q9wA9QJBMz0LbQJL3WIuWEl71nc1jAEDXCGNCU1/xFP
o5zlc4GHw+BZXCI76aT5McHjOKRW3EfFs1mhcQQMV3WPVwMAtZ60W41oXe2A7ZXVkM2iZNx3R2qx
gor66GyEssbS/i7F/rRyd/G2vVtJ0pmXaI5DeWz7dDCze75YJ7h3XAJkqkAzitr7pVtwZJa5ec+7
vGjYNmuyfri/3/0SpsJaTdIYGo1xsa7qmmx+XPiplgOexpUcQ4hKZWqZRsqQ25qrvjJg/Pno4Taz
KYWomb5uAp5C1Tmlxqvy+lxUNAfzhzRgPOn6gH1K2zFiIRMKMQhsWqnUd27ngV9AEqrv3/JCMDAr
hzHNiVcJ4uOCnFTcHVc3bOz2C1lXt4OtLtVLRPNF1OwOGNgqNxLiwaF7i0Km9s3/Jp9TeB0Tjo9k
VPl00AmUIKigx6AQi0/BP4jZRJ/rtZhIqIHKWxh8FSDhtHCyIfSHP+cOx7RF02HITWxeu3Ho8I5a
DAZ972QnykYxnJ1PsBaXOuOqOHIocrPW9H2rVdDST73luVmhhmsj5/L3KBq80SJ+PS2c5NpJ9igZ
RLHchLhyRiX7LJey2w2aU1A3cAJAyqzXjSYpquvvrrCvcsHBCe8kGmFlne1NlPRymVi3eZCo4ZIO
j2YSFnQZseDl4VJvwRPrneTejzKlTqjsMJPh6sItWq+E2fkaRmVQW4jM4wmixxYDJZtyx7IzkNkO
n6tHFOBGrNND3Czetrc9/gakuz/3nCvjx5vPN4BQy3cWiUhCPhlDGxpGhpN6EFwAaiZfdHFw7ea8
gTFX6BpruPodYO1fLiFkYyHQU7XgwGqpKs63Mhkwn4Z60GcOBttZCHISc5EEtsqhnQgPkS9ULsBI
NIfEo5t/P5bsM+aHcROiOhPhWRLS4jWHu+v3T5Loc/YMnMZsfWhKqGIm+zqps0XcNpetFz5lUzYA
XlZOUJOECAAQekU4a998SaIhREg7HOM8FpG1FIVrb8Yz69Il48wAwh0WwQbQSg4lVzcCdwYKYiUh
hRQDVZJcnGGQfOzNB+PaQOWZYAoYXto8k7ubKYrVg/4i6J+Mc6vtB71pWS6/NcrvKsMmtBo1O/l+
L9XpYwd75JfNwBUAizry3pjoAeviMmPXqPwWl7PdBIhARWMZzFzCxyWqXS6SQKGvTd4TlulxC23d
H7tuLXWBTK4sl1Hwhse+wK3OzEOhim3DczRYIKRZkIfwmrxO+erfrunjCdZgwM8e9TigemAPqOpa
RDly5u7uRziQvmLMfsDah+nG3O1RKzeQDLkYBTohus4v02g6i1vtehXFwxVHb0tIY6w68j7GID5P
vTKN10AdFZIaQepSvFVrlXYYP6GnIYDNq2VTQuhr9XBShRTHu5ZLLaEiNQJYLdqY6dM4eFnlZ02V
I94YvvC6OL4WGAe/y7bUPbK7TrKXIDYIDJ4mWHnAuEc1Uh+v6O/3kmrd5U6N45eA0FPw1BUKfFCE
vMVDwu7XATiUqqFCImkWNpTgJ9t7UyQjICS9qUQY2VZPnhWg1UKG/1mKo1ZaEnCyFPIs/+dQMNuM
jQMjXZFFe0Cr+vYyTL4FbwgJag3fCBpsoCgUBltHA7BlUU++snwdrLwUHySyoZ33SKjPLJvL/Mu6
Fimx3ZyaCeAyz89HHEYxJMIj+K8iBR8K82AzJqlwy9RFX7bJ6JR3IuFf4siqZRHSTgwDwa5dvXeS
dEdiaEmnLfvkYR+f5tIib0nXZtVGXdW2SXDaAPuyTThIzHXGbn1S0lxQGRGr1/5/V6ZE0old0Wus
6XUGAjCNMwgXoBRaqqRVZO9vuhDCKCpZB6RN+bUG7B54GqQD2qUz14EjCLbSvnJ0Mw3wP1IqREWq
Iw4pvzOe+zat9jS7GL8DL7s43n2GzPqvGszteHRmmlwT9HsTIK8Ipass21t6EYXkhHb3+NRnPhTE
jh0wU5RYfw6jIhtOIj8qrclWLwMQ3c9PvmTKXrN2fe5pHdk8l820IKtmyQNvRACQiW4kgl3B9mHt
NmKXPh4YbJW+47HQ9qc2AkkqufLfuWif/vzwQF/LA0E9wGmafKioEO75RkLQf0+7isloW5Ylxgju
G3q0laJEPKhlUMPtUfgNY2fmMl9G8trGxE4ExfYkdSXZz2hYKiNq8q75Omct/vdGZfqb7cVcEzyi
LK8ccRfQtSFdHn0AtE3eYxu5WYHTeNW65OR+uD+9pcivEYS+bZIHMfJGkM1T024wDutt2iHXYGFJ
AfGtzP/As9/8TJ2YX/kFoa0ofyEKm0FhFygwo/Zq1VE/KopDT69GQQZskZ+IZBiGT5JRgU568Dp3
mPYXTbnU1KQ5garLqRbT9gbklv97/ChLypWPkqJUnnW26adH799sFNd9ZGlleFKNdN0yVMEpgQ+N
6uG6jYuJQgs0CJsSFIfuGDLPN8WbBoCgtx0KivWChlbS4WcEq5NUVJJMlLVSFUbPwEBkB+r5B+OV
Lg9uJ8QK6iweQ9ptopBxjCRAm/a8p4Q/LRdzSdK0pWBG1i8gOSSYtSgtBZELyWpem8UmT9SNkcCG
blcMO/DGO4EV/52q5alkLGEG2wUeFUVWXYCvOus1zo26iYmoEZVTW0tmIHtVy+qxzqb3UY6Ce8ZV
YXSl1CP7UCxQo+qrL1ZEboPZtaPI5ZhZDeZVTxvPlIRR9T1JpIEwCRFd+6DXl+y9GCsN0ha+h7Yn
aT856Z7CnXywu+cDJGwz3ffxzU0SjwkVgsh+o59VN2C5XKiL6zoFBQZpttzKHm/Dxt4a9Q1/rAfr
u82wkFGb1y7AZlQw2YQEHpw70G3SFyxHZ5htYhM4aK5RoWppt42GvCIHsPU2dQcj7zL5K/8xFNot
SG3COq+pN9amMOW5g17+n3LnDg0l+ElKGcYpbd96b85KOuRsaBWFJ2vtYwWyNnyjrMZCWp1d0IsV
fpyIGiBSPdV7/2+12lO8mvHO+xORT6VY+ekTT4+yQPiIMzvtUecym1YL5DFYfK/2f39YrTOQKVyM
s+LFwYWveV2BsvsnS5C+Xd743Ox97Jw7RgHBY84y+aTBF3wC6TYN5+y3IUCrbaDnj6VOz6+5K6Rt
virZqH9LjBEAibqKtJMJhAoFEgOjfwfceUwpbi19glsDOkwFvDhB7zq9B+yCG2wHQWWQpBFcwmI4
cR1ux/6DHw/GHf/l7CYjn76yrzSfmYSvhXXCbGG4HcvARKIQTYb3GyqMraYvoUc1Kwax9i34YBxV
xX0zPkA6Rj1/uFY7P/0fuel3mGWPKA8hrMQ1fgti8YFs7BCH9ByrEy1ReMwrSGPIbUzx6xGtY5j1
Jl3MXKequJ1FK1b7YVOP3FSQDbA/V4Q043i35mOw58ZWr/q+yli6tYqyP68ELbV9hFKj+ADkFfAV
/wlv+syzsvetfSzeLQMK3lWMwlAFBNRSXu0hhksShIrnwRlFxseiaQiCRnexbWyJMoebcuHPr+k5
Y5Js5y36zd80hZoiugc87C4NMFiw7u8EB6ZfWUfXO3MJQZBsP65UF7V2GhrlOo8+V8tY7uExd51L
GhywCkTPJTkT2vmFs3KZnuh+mk4+ux6bQ3aqBwgYbRCjDsfMUTtoibtaVmFxbvuu0sW0xR0HOJUM
NoWKKb/KYdkv0ZC6YU5NL7gIp5C4vtbf5k06tSDgQO4RAp+T4y0FTwlV1+4wu8ILKk1tuZDUoevN
O+txhPr3X/0+9R+0o9PnLWW85HEhj14Ik3tSjGqE+JYIuOSxhBNTabKf+UPCEJH/Oeg0mvYWHoh6
A4lfBC8MwC62ae8SJSd8KMC77qA7PRFCzeyoF5c6zL253KYDEQE7puqowlm+lS6n+nY7tOoMUcvZ
WDXu6Tou3M9mZDd5xskz8sisdNWHppfqKLdm33se26VLelVxRsuVtIXZCfwhc8maZ2WNqZ8GSPO8
0CbEs4l90IvXsxA+hWBS5tBHA3raLSXk0Wztr6oF9mt/0keWnK6Tr1V2cB05Gd4WCxug8mF7wfBM
zVSYXcjdknNIgyOsFjlCp4a1wycB08mlpEjoBW4T3YOO16HGWKkSi2FFrCPE5Bw3fQ8scC4TXQ3e
UmfCZX5l4mIp3bijaRRJkp1DWwTWPNBxxlNHrIZ7a0y/DPCZFNEyY7vT6LAapHEE7sz5ck9ihPHm
bXXhLrijbzo5nmPMmIFc4MB+5S4abQbCSdTj+d+lMsRNM7HpuFL4k0Gf0ElWVbkkjgPMlrzspy/L
Jo8CsfLa4jzZMnZilgKLBY7k2k5osCjWZ5sD5aHGwEnoHdD9koseY5thvehfsQIh6WKVQCaOoVSp
mVyLpKtxv3hvqlpE0hkefGDlCpGWsMWyj0lXG0/8n36snT8L5aHmEssXZowF8mph4IJOt3sK/on8
WOHuYIWCsZjf57QcPGtjmfxb3ozzMkKr668v6IcMHCL5aLO6YQqOOHsjpu2QUPVYSIt4CfA0f0lP
ONDv8GZaaEJt9xTLdm9hCUKMLXv6TvgHY7fFq3kJ5zeKwhrPCBvaR6ExdSZQwhoLEskLakNNpSY3
UOP1UAsF1uemIXbRBuYBBwJl7dKYNpWnFuxv3Lx7ryVUj04a7nHnkUMM+ec7FD/FmOpsJGYQdFRZ
8Xacl0rP+TG1c780eo2m1liCMrWltHxU1gkez2bxg7cxD+eqUFIOT08DzJ6fL2L+wmXU3I/IiYjU
0Ywf7m/Q9wHfNzkcm9hqhRKkR4ZU5IdRRvvx+nwgG3W4sXLsNTINWW0lmomZAYCWzJo6PbWmeNXM
8zOArvlZNBAPTIm+Vp3qhNI/1OYgUeKEyLlh6dFS8+AsYhDKTAkHb6IrUUrSQC6Uc0foXKcaQP27
SD/z9HESUW78lxpigzWnOnCMysZbZMhJGcBTn4vNy5SpRaB4tBcXcJuh74uMu6SjNmtFrRPqURn+
SVvCMVQuX4aNqM56Z8xM8Mxy3mJyF5F9yNn/QRicG4QLgGUUDuCxzb4l2yIrd+GwtQB9dRuSjFyj
0Y7Y/vOUKTTkRpyVYhsDHGoxVvIaB07KuCyQgb8wi/2jq2mBoRp0TwNSZ+wDVUtJBPqfdFpeuJy0
84yLQ/YJYKfywPXwmeZMnefxYxyD5sjMbIcbfrUXH9pbq+f+BFMBfD9FI/KKlP8/qkUl61MgNuKs
yGQ4wirGLlzY2OViYcQE/lr6Kg3TsKLMMll86RWiUNF0/Xx/NUXsiiq1ghVW1ocMCVnNnHpvYHSz
ZCVskuZRkfx3iFeRlk9EPOyKKemDsTdZr1a0Sub43eOIfP/3doflPksdeeeQjVpUWmpHEkNVPrdG
E7VDKPcfyHWx1OeNMOC8JlXFzWvV2MMzYQhLFDW8BCBKG8pxEazMC6ugmcZYDNGubqurRo9SZZ9C
kaGqIHeaDVIBSa0QZ8zaBd8pLFYhGzfjAKUymr3CnT6TfSPrbFg55qSAo+7xPqai/DGlGFKCve9W
RgK2MCv41+xXIRNbibeJeOcmngPnKSx7+//Zk1yptJSgohI7+oOI/ITu2n0TMY1YgGfm3lgf546Z
dE4BwlbyJkH56xdNUPWepQF+4YQe9aQ1vzslRqqnBphIN3XourHmxGk56hVBtEYjEAhlmewZJVOt
TVxZfbow8AmztUfV7O0qVPw03Z56HKb3xIa7AdvuuoXqM4tbtOFUL/k7tRv/qXya+KxJycQbxwes
GdW9ZAkRP+85ZhN0qKGsLLqJtkxiVEG5WRhZjG70h91QH5HUinRdXciQhWgnyj8vXrM2un7D0kKD
Gi4FnSSkam17jvneelGlIK+zL6/knmtY4UAlzvwqnX0loH8eMHP+gxwK4TVNw9R1NL9brr3Ck0MW
KpWvlC0fNdnsyMXP3iJdpuMMsHBsuulUs9lyNG6t8yDtQn/fZ5thGKkc8rEgp8xM1pw04/jXZry8
IAc77MGRGKZRtgoPJGdW635lRKA03+xtB0qpTKTJm0r+D1y06AvU1C40RflGLGblbUHvXsqVyrl1
yQdrSRUDiFgQyAS8nQUatNPLN3Zz5E/0TjisMAkjBM6GLNOa9caAOKHTJjthSXLw733WxQqxJdQC
dfWFvwKQ8YBZcoJYjAasrzXpJwp9Ia6rhTSZ0PTbrYwEasYkQtLS0lKbRRMkRWNcihV+1VtcZckX
pxOtWpe4xpDZ9kvNly+nFk4vrQ4W54K8LFZba38rVpxplkV5ZOyhVQjsX8rSfTBsuJFw/wIpwNqH
+7JKY8460kpeeUiFaHGIJ+S2PwPnX5N4K9dnFZN5rguK/viRTYLAomWOJHrgLMchBQBpVNkREUuC
P8o7/JBEb7+kjsZJBEhl1rX668bFVOTce/oVijx6HMlyRstN8/xUQK9Lj1JkQP/3zbwdHYrtOtpB
TV4zk0wfQmL6ckwL8/xqaTq+wvcNeZbmH0Laiu1Vl5INK0pH/QrjqY/EXsc5iFQNmpRkNdow9bi6
ejdwE61mFCvBPOJFdnd0Fx1iDfK/w5dFcMuj4WBGwMGz98XqTB50X7/zF7gzm22xUTBF8E/0tgUq
+ZQV8GPLm2k4fnaNCmezGzP7X9xe5f7I1Ygzfv0v2iA+MHztNpuyAp1/axbgY5DstBPbvRWfxpCb
EtSUZwYAEUxcGAkrdCvhEFpaV++wDYAxJEHF65IFr9rno1jugdKGueF/NidVzVOsXsbm/8tubHYq
ePOref33yo2/SLOogAHyk/MnQc86V5MDY/d4veWTBGMhT0iIZQicYNoZ/Byn+ZTU7uWRZSB9tdmQ
EyrjnbySTrT4mzhq73MmfGjZZdCMW1QLdFzaqVItzOyEgOtQkdSWRGKjjWfa13Z0e8TcKtGXf9Kw
paf3fMtfEzTTtV2jGuaPXv9DepF0Z3qugKC3LNpg4UMXRU2PbZqStIHxmmRRCCps/MGHfo6N9vJ8
d4b/dqnWZ+tzVztKw1wZf1P39iyv8fzoCND1iYW5lDsWYz8VEjHWgUOR8vkjE6pAtKOBqxhMbcQw
QyQLp+dk6yIhlDCHNUc35/RQ89IEiFAtY17WiXSRrxJ/6w0mLfB/Oao7314NI0ljmkuAr2kZQzgX
2emxi7R/76PDvg9AFa3LCKzFWuqwiMbuSdK41ZjfvPytPbmkN2qymbAI3kunI6TGlHls5z4m+v30
mIMxvwihpL7SeAOBLIDG98bObLvl7CdSDeoMzr+l5y3z2Jq7aqwQ78GCha+mxmOOBFeZNUS9JB2a
TeUPs7SetVBrkkjiu+KI1XJqqOOjtHkMJiLRNYsCT8b1zlUYQJ25GvhSqZOeWf8QU+ZoyRheaFsL
kHKM9Fx2tpmcxVEzqaWnHbgI9LJWsc0ElsqRqYOVhrly/szyB8mPeRvm8dtdgbGmSZPOiP7J39lf
gY9hnkiSjWBstZYgF4x71i0W2Xpckp3EFYJwoVmYwUFNvBm9gxfUfzGqpDSC2HjpqW1pXVNirwTz
fr4kQ7yg4GonAcI/QDG3v+ROd/nGAuFs964p1uluiulVOTwyIQOp8Sdh1rtjPsgiuZM8Lep+EGFQ
Js++bsFWFYCh7XSvu7FZazJ8cr3YEAUGZG3+2fQFdP3O8X7Xr5ad9skqyW0nPR8o9UFrDL+zz84M
vMdIRK0//70RuuhlH8uMzeSuMQ1ZjU6yo3T4nZiTMAAU9Gvx4KNkvpc0TeDgqsnj4Nt+1dDO2YeG
yLtqGNsPw/rGPDQagDb9lU0HaF/49H3vd4A/4k0Rih/H6M3db+NiqWWEPFtLAW5n7O9dLQAwQYJI
8ATSj0EjMCXWUN4OQusq/xfqNvxv5rTuK58bMupqPIJOpyR7HhD6nz1LWaUTvBcrfQg6slpDSHi0
OjbzZHruQmAuH/13veLu6JbH5UA/8LKW03Tq4tID6mwyDicHFhBVkF0/4cCAnJnwO2HN+pZaOCn+
G0H0dYTpQkritnevkdGSPlW8cJQDo/KURBPgFq+ohixiOH1v5C13JO5HKomSyvTpbaKa8WZTG9B0
Wyv8hwi+kvfywNLayASstl11pDVEgZ3ARiLlND+/Kmv3PCFzpcDS5+CNyAcou/re/spbtLSgTn7N
pCyXN9mZvBUzsdOuu0OvIachJY/o0aAvfh2OrMuLSRx/+Grb1e3gSwGAEYaF7YY12FuRLnbENi/t
dCFbA8vUlHJmjXmseZrs3+h0RuEaDQ1LDgQmciGPux8TTbs9W1k66A/ebGr6otH7vcVqla21H2WS
hn69rH/fuU9x+BC+L3wWaGFnQsI4lxlyXS0Xaqp5r/G/TaOdcYZ+1yiP6uwufg7LcDKu0AyKBZ/R
E8atwDcIPRwj972OEpN2cChUdHHCopnu7BKGBCxO34xvI0WN8IjGtXNerPRtBAjnsjJi1pNyaNCA
x2q4ijjmJbNppeTc8hwGPqspovVY2mapKHxDnOHworJlCVDsQcYyrL/pkDGwtz1Gb0jnjlLHT8cB
ZwLGlVO7uBOJzACRBRfuCUztoTAJFckAtaWIAbLA6xpU/GAob2C+hYzm57a/Xg+g1XRvawlOH7jF
noMcUDvTtuNicCBE/bXpoGwzHcjeo7VzFG7SEsMIfZ+r1iMka3EArUlW1g+eBjU8LLHkjjPdygSV
PT9t0ZfPafU0K2Y7M3T2jud53wWlutBrZ/8QD1yhEmK78sv2XuI+xaJ1JU8wBoNKmVpkliIlTWX2
YlBFpcPt8jta7/8hVf4Nt70Ik82scJ+xTY3kcOgu5DdDhSZ5oV15CDWYYnaovFg6KCjeYHp4ym0h
0mMKxpQYvar1gMFgNH+F3RYlWiAXkAIqg6EgLVTK8Wp9NcC6STZGFk9lba6euMnk/crSEnSXGcAJ
PVlpqccgAsvUrycNlK2RmEuTSvhv7364oRLFJ6k+JvhKgw4M46+wvxD9130ui+Yll4prDBv3wfkR
5PYlH8h6nl4ZBhkKgoR8LlEu/JpZyTOBQfDICA1cZWkFjMJ2ShHdXe4Y2DqL0tX4NB+f6h/xjyLG
HWc1oa235SE/4twrPGBUslLS5bPsuStnPhu+h9uVDMQBgOKIEv2YtIlmfbwQ2SxpMFi57H+/2tth
Ai49N/rOGzedjail1r4DGX8chJntgfuCUpD+PKpQzqJc9g4kO8tS2jztefnALyA6/RNGbwtnLb4b
VS/nB9Om7/g5Xo2/o92QtFuqRdoxBWPt4hiVY9HQKiOzZPeOCU9UQcvDqr0ns6+zY5DjV0d4UYI7
uYN6+mqkcY6P85CDXigi2xErfDYBmwmSMkvt8IaSLwJzPDAQrHNx2NOeO2g9wSymejH0EboPTJMx
2o1yykcqxxq74Ejowy43I0SiOO8Z1gYNXe/euLqXsNC+VszQx6tGf+8ULayv6tMDk5LBZKc53C6h
RJZ7IoCCknxuS19hT+n5r8ukIhf5N/PIh+26zURYbWW0xk4JBxIgHzH8FRkdueWhgHj0nb5Hujji
BCEA03acoXYp5JK8oke16G/eOhpl/NlkUq0MFmu7vYRtZUOSCCDrx6d/zSXCPmWXMHwyD1gG6FSK
0I9WudhCkVClH48GoeeVWmCcrZvMYp9kv20Z5gluoRJIE5/mceJLxQgkl+CmJqsiXrwKqF9C8uyH
gnTwEqPe5Ndyj5HwFgepW2D0piUYppZsPxMtWVuTxMeqQKz5xOFm9XwXo5PZCGgfvIVJTVTQZSgv
J/wo6170LTgh7WN56qEixjY4kTZUGXVwVp1Tt3oQiEaE8tlswF0n/aMEpmLVxBXVtBGSzS9LpgcR
bOz+VX/EZfHH3OvJX0ZsXU3g0hWVtuoSG4Agx1NUrEHt/iR0tFuTpZuPK9WVos2KLt2mFoBpRb8M
GTOWn6RwYB8agYNbiUdPBkNCqVxQHMJN8vr9KVZil+1AFj8DyfxYu0G6iDYWNitB1ZO78z+6nFou
kNwANGi1dI1BYWsMEXte21dVR77btr5prrTPOpcKHhA7fvQ08uRfhoGl2N87j4DHAqZGP0EZwwvh
EJ+ndAUCsLId3F2l4xiDheIoeVHX1htajURG8R+qP9pc3OCK2qA/FGyXYibqyfjKg7zToheu3i0F
r9RQ770/ODs7VifOos6MGPVPVEIAlASrWPx+a4sTeRW6+RBYn/py0rlmVKL0dONHwQt1shC+eNY7
Dw0U6EFF+gOoTZ1rGhFmWwC8K9z/Inx65vCjrIL/kDv8I6Tbbi6UzJoTZtHBgdyUpT9hHvZHBc1t
Je8FDy4h6Rb/C4lgM5LnfcIYT+vb/HWieDwYzXN8iDRxhJdViCYzapG6Kp/euTH2o3+W5HhUjLSx
arx5XPXFItTXHdWH5Czsfv+bNez9um5YZh7O2cXNIwwfyFK86RG+kFa3CXJr0xq245lzgOF32IJl
vtgPeEMibD+upREg/1Y1KbIXddxlA0eRr/DOzxl8xXSvZC5VcAQa7OVTuYsS5j/WURGm7+CNuT4N
mTaAfvzzAw0bpbJ86d2Gz8fnYuSbBQRU41WacyuSPhi9adoEgGg2DAwDh6uwdej234JEubeGNfoF
NB0CL94qlzqQI5gxsKkK0St+D56PVjbku2zwpkmfZ0MKDZbfjULXF/2PGkYD68VaxVTqwBiaKcfF
1NLslHBsuRNYjcxtn9njEzSFER6OB4YpLjVe6FSqcP5r1JMkgQ9kuhv2XHotTgE2bFMpiryNKMes
uIPRZVJWUzYzKIYYz8Y/1ar+A6bO6qhq41O0NCdJv455Yu3INo+DbmNVrnP0FT4vg1v/DoWalDTJ
EYWGA5VmNcq3stvx4zCjrFkUSBJPOPpCmRZt9j5yEyEMO8rf9ZbIz2MIx7R/CzG4alSwZ69+ZXCv
9lsa0BEXRo0SGLQ1GqApzESRrzA26kaqpHI0EExmFN27xeBwI7pgtUb1C4pfk1YUlfShGjKSt+sl
IJ9+/p5bsp3Rzg1bKSAF70fsJDUvQYHDewXJulkD0JWPYil4WZJUPTfCossVBAjdcqZ1nocoBTS7
f4iiHjnJrRjyo8wn5J/G63OR4qx2NqEbhU3Sf+QgTPNh++X5boivpEt1wpdt1mV87jlGRrsYDctt
DmQsoQKWsr+NeYEvQ3lgAnb83t+9adNvQixeCZub3xcIHMLfbpFPrCxo1QWCXfDTBeUD1RsjfuiX
moMWILaGQthfFpPhvkJpQidHUOaWyhjqXCeCz4jYDvXkL0L6q1wmOSFGdeM2zA+ogvv974HwldKZ
GSN39QhOgmGATXCASgVDY6cSmgJEwYr9otE33ok+aAhUc36bqYr1Vk2mlUYOdw8XcuoC22USskRN
1opJ6glhMqWJV9SzOOC2Nob+/+/LNjVIKdhwJVwRo7qGjhfISqrtxXqK/3UAoopE+zNl5xip376b
t3RqWyMjKpNXfM4i8U3gHzcbiRSvxt20lkhNoqd3Ez0xZxTQpMDmDgk+PnINsfqDGdbnB/IhUXF6
bpy3x5cELCHDH9QBX16OqbNOp0wMUtnvTAdo9kIEcnmkBOjRIlXT7sdOH6GelYVGeWC9XeIJOF39
mbiNF8S2uJ4NlRSK41nEj6j5T3WllgYDtgqRcwRJlKexd9/u1JoHCFhDeWGIhj9htXnKB6oKnTJK
Be6EmY3OVod+k5fbKM9K46Dv4f4hOF5O0dFOP0t+r5FnWYr1UTrmI62QNAzjctU/mojHcR570XPU
HkdDbSjqzUQ7HyGVvps8o9V2D8rGX+Fe3ZywlzlJAgJIotlrTiY3vIF2++EiHEjLMQHMrCTTUT9O
Imr3pG6H3OPFi2sxqIrJ9BB9sNTFGabOG0e8MS23kMF0Cl6pycb/qydCT3n+gItlLzxNZFE4RU4z
5bGANt8Ojgaw/d5rwtt82y5093o+TcghDgn/igmYA3OfHIduP4sbvMzXg9Okn5jzPX0wmoPlX7KD
8yqTyeOgj+GfihFDGXtEbbyHxOTI8p/hWotuixeDDgHlcz7QxSPp4cbM8XWxCsA+7eXjSQI1BZd/
dKVpBB5Ry0ry25GgmAI5yrJdG4b7xWjdIA5B808AXXTgvfBWZG6IBQWitwFDor9HqhNrx2dfbxcC
Lm9Qq52moUsVC+T6FUeUG+uK/fNNvuLtXLK1GGg6l0zRHGhlLPbzRyk8Nu5Af7WYrfhP0B83jhhR
4kJvjD/7ju3FBXu8Gko7kzNOQDbDwD4hw+2xj8ujnGd+EqW+vxLC/BxzAdVumBgL4ccqhxRn92+w
bDltkjDW0SSLfKpRJwa9gsOnmakF7Wbum5wQXyACZBC4E+QOdLf5ZcDtrfGNXSWICKGAhSySJoGT
NaXPCE3E0c9nW/WjNkvNcIw7UvyxOA7tnM9qA42dKizUN0EDwqG8CjY7a/pYm9cJjogiv1l/2O8Y
6lCJpX3f/3FWDuywaFyRbfvwbTQUEyV6TKuDI8t3kJkWWhlWcc0/6WYMv6JzOcBFSQn9OtafOik1
O5kS4Md2aeX8dLIJ52aka3HkqZVYOoX9w9iB0PhHaRl5ZIftyuhiIwi9KpPGIr5pZ8yffbUNY2iD
JXqG0c6oJ7eJcca1KNzIo1980MNO5cZR/VUSs1V5O4n6PJGZURwuQ7avs8GI1A5ev9W/KBepjwXS
kLNB+YqlYEsyaoCD3pDST6OgZTnK0VAnoCXxkeSvSnJchZplPJO5ZOj5ZTOaoiCoKs5tiCmnFjpy
lbGWmI84AyU8jcegSzuhU4wwmVNv0SeVAUnleGuEZNCk1F2Nxk4G6b/lSm2uRcl7RCw6mohZ/M1d
3XUC5GBiFSlLcv7KW2AwcKl1p50iurS2S4ELPT03GjSQ7xEiOtvcaMqlEhZ/AUXU3kaCRoE7234Q
w4PXeNqKhdN4HfePQU71Hh03sfM/QvH0akBHAaY7wwLepv48HcKVrfq513WugX9KrMY8APvoMILv
u/8AgzrjUuYTC2rPzl/gVqIsCmO9xOOOxoGX3ehtRWETgaJXfl/I8JgvT1ILFYUo5cURsnbjRyHq
fIB3XjSAoau7vKTvLyUdkQ1xo3N8FMbFEtt5aukPrYl1QEcQ+jQwWXpzM8XKt5tGtxCb/Pe7JLfe
TYuZn6f0lpafW+1YDge56iusSOJoLgo2mD14W6UCLrZr+Cduxz7ryTiN312RyntLtwMD9c7wr/9Q
5dinQeGnYPlO4hlMamuILvKYSEwvsk9gO54osQsRxiAGKR4pkhk50Y+xOE028fwOIyNURS2Lw5nV
/fj90IHZuyjt0UkQg/ynmg6mwXBZPAp4Wf8zG4bjnHTzc+L68Uc7mWU2nvjv1TttjEcnsco/Bepf
jVQMIyyPtai0ao29y7aAjF8GxiVA3emaSnN6DpkjXGWEuw9g7T9leakUxGzHa3JRKufN/WfOwdcV
eWLdZqBMjpF7VxRcHUKRNIcgas2U4OvJB8zKB6nrJIv5Bfpf/GXKhE5EanLhB3Sr2qWVFIs9Op4v
M42wLX64tiAljEWPIctOyAMC+iLghZvasOAvY2YInfuXHFwfFLuPDKmyGssffVORPSvMJkjPOnSt
c8QSPOYzQM5icWaTZO9YfH8KQqKwg1TyFP1QAQsGlF14+9G/l3pcOxVpSp/sWSWoj12HaCvScIvd
lYqqHFNixxeqK8XeqriiqcEJ+xkMMd30avq0hj8mLMKILW2w8n3pDdMV277wxeWLPEEu2fdBjhUA
e5v7QZ2cdBuU/12dfXw17Ctqap+Oi7yLW51ys25Re3Clf5qxGzkZHcvpfW/KoTQrGDlIYyxUGZfQ
AbJfmHiERnQe99nT6md8Rd1SSV24SyUhuXFkesxqnY4TcOLfZi1pRTbcSgAXqzWfYELpYD1FdxIr
RGVmLfP4ilbAZGxx+nyyQbSFa4TUDkqPwnM58pKnkjdYpTirVFQbFmkFTo53QUOsY87zPkjON7/+
OZWqluUKHRACxKrG3Iu+utkfvSG52+CB/PGLRoW0ZhY6D9VjhgocOkPo+Tyve3xl27soKz9za74T
UUpE57KlGadXQgrIb4uVyQNt3whQLMEe9vBv3pXzPVab8QfgZ0d5yTg/4wrWXvh1ZnoWXfTpAYPI
bjHFxzHqebKKnFTSKXmEGZiKqB/lsVQZ6xCgsiqHjwFuOPoCqskRv2a3dlAv6ioC8sm/TBLxjIlZ
vLVxLNsKDmp0CQ53ycgub3oFIjjT7mfOAv/6QJHLV4HBSW40F5KENabMyaO3v7v97PvOctB7dywp
SOl+pjBCmch7skJ11GAQgSTb3UejMSu9O8SSL2U+LZcYNTFv4Q27nLD6qiFppe67I9p3qsnrwW+7
CZrObCRxqW7iKYhdo+qwmO1i93Q0Zb/mz092fupgoe9kgebqh8Bolin/WCMy20xAyZXFP6EDcFIE
pxgzLQEZ5ZbhU+WkWVoXKMpuJaHgUcbM6iGUxnQLBgus3F6K+icL7HhdBHTTgRPnbvgOoTLrVA/E
yzwPPz62Zb4F6Qu8YfYpql0gm0Sx72AhR3Aw8HnnnFJ5e2YUYFtU7HuPTB9+FDsnwIJIT590Gu3c
g366JXPmDpwYNIdnYM9HpRQ9t1z+EUeN5JCXZZJEwwIoVpq69GZjNugD9S4BYSlzRtE0tlO27Zs1
LhDh8y/KbOHDKXUWfSWOsJ4cmnn2kvISoumZZ8UEhiceP38DDJ8pxuzGAX0m4PM2HL93jl4J9+1b
pos4mSzsvS9ywjhMQCaDVUtLpUqV+Hh97g2KiS7Pce4S1WOTgeySFypbXxoAu+qEAQDblv9jKD27
buiqWPay9qS997R3p7BqL/rOa+lW67cxt5+Mz7lMDlXyA8KghKwsCZQotYnMy8qR/KK6c+0QSUje
cTjMuG55Cj2gR3X9j8Z46Ul35/CNquYR6ziJq4tzHsEkP5pw/gOmCUsGL7CEqB4n0JshNTG5zZeX
GgyHDMRlpBe2qGKlZwZkVeKh5D8r//eSaEn2Trz8ElKCo4kxibkIqAKCHbn8vQaDbh+gXZHe5WCP
IzIPshGUdpexw1QTzl/7fSCni/2EuviHcM/liGuf4SGeqzk1iQobGKRQiBh6wj05jNdOG6XoAJCT
ldtUawwyBbAm3lYrh19ENapzCBAA+RV1bvID9AGIIW3+RgZK1zdIGJwXScFYO4yZ8p9L0Pcqp3Dx
g4Z2tF/Y0Cdpi+qj/2C/v7kHPP9fYQxt1huj9fkD0REM2/7Ces7AVSX8SWo1QjEAUgUUpvBVOir4
ScN0uhtFaTku+imeGqO2anZMo66n+Ar2witwcNWZNkaIPeI59vbrh12Mf1DPcfO4MLz5KFwMhlE9
D8M6fd07/DXcQ9FKcmvNmy33vlTcxBOcHYDMG/Ys1m0aNHQeXBxLo3X6Ackb55gAiesLYg/qt5OU
y+Pta/rvkNoN4FNLGV9xp9VPhmRl+vmAwAq4OErgDl4diYXIidLvVt9cXCaNPtErI4FvBAKtXtiH
ucoHYylDXOuxOsqWUzgNxJxhyx2EM8P8pmrO55k8EcJXBvlXO8FrTErkCNiHxHaGrUv/a9F05nTC
2PLBHKfjFOvPZBy8V2RxoOFabGvMk/YBiKFtq4q3y1lyzp8MMDeuk8S5igBKf+IdAz/DIMEL4BVt
sqwzkBS+cvLLLgc7QjLIXhxnOk1MKZ8iJi746kCfkEcbIo5FxnnKBV7/WZUm8B9uVbG5ssQ66RrV
/mw3t05y+3bk/Ut1xvzYOS8ppqeKGfsDNOdiSLPEHMyR+ZHdxkEWVtTVmgK/txrIps+WQfbOTjP3
6YGLdIy33oGMtSWf1FDbWxEbtmGTc+u+cONiYxqkRuxIT0W//L9nU8RY+pqN7pt+dHnFkOUw5Pn/
R9Y/1OZLCwnJy0rimM4ARYiXWtJOSaXa3urG3hcJCI3DpT9GSDmpQpDioJyft/AglgJrzEWKE/2r
AzW0p/XDAH0O7SfedBkOc95ORWccZCB3fRXoa6amo0w8BBGqR57Lhaag5QBoFFJNZi24ywqos2aS
qju3QWA8uLfIsx3lGixUAMbQNQQmlleWpTbyQD9Fgo+8l2VNOibdmOLrRdNMZsIAbdhZgVjPADb+
k+GFGlQo540kF8niUwAHwqOAuniRsayT64Y1TEzlT0N7f4PfdFZEVSfSWfjwIiUVBvIGefOK35M/
lZtXFinM3VZFtQI3ScwjrJ61rx7puh/HMSfGYTipJFmvaHGAqNx0M878SwhOpAHBckPmOc73Pjw2
sXsNqEsCr/I5Q7Heg6wz/lrFnib5cWN3eTNVkIAkQwmSd1fHXHhkDyTnNrrOsns4LZszlAdqBdmY
r+QuohRCPpUJ0IWAMoAG/4IRNed8d0knucbDxE60RYocbFE6LGWzSiosAlnyQiPc5t2u83vQHsqF
wKNKP+r72mj+1uYJFLI37qz5fVimsdJ3j3TuneIRdZyC164P9gOmX7s7q5h1VDz6XMcDMk3/LRBm
hfOEDRZKeGyweZ8wFnhOxuDSaWeSE9Mbd5wn2qlNKt8BP1la3wh7ZS6O36SALbtUtXstkzc0+4Lz
r7iaU9neb9nbJCsbKnTSiuolpnyWAHNrYEgcqXbrFb0Yo1iUzrqc8DWlMfakRPJmqwoM7f58bkQf
4HyVNfHU2WQJwCexUi4sCvwB7RidSzaOremihorfuhrYS9m6ZkDnfly8x4xJPtIOrFWoJaxhxEun
GGEMcgdkv0QST9COCjSigxStTWlnvhXMgt7kwA/FCfHBrGLBNXF7zNRRAIdiDDV6XE4tRMv8Trtv
FTJF/izuQdFatsxvRDPUnBCo3FlZX/4PmPHXOxFdEAnMJri7QsqJ64LqbPFZTSK6Wi8UT6X8H1lu
0eY6vHHXmIAWb0opnHoy8pJDxYs446CEO3ut7USv45a0T5LfHWbgi6yKZBJhOAaonyQOCwYLlAgk
qJwnvwoQenjkW+0NUYd4LQ01RBy9Hx5kjtvsSviN5DTearWn2uwiar0t33tlGH1c5Es5v1y8J75O
cX8Xe2lZhok+4n0a7kSit0p4VQJvVbE1op8J3QamEHXxOhjLSWuJ5S0i+33vJsM37MnvVHmCUW/d
T8At/v4I2L+6g9eGzgrCMNpjrw9IWBGLUhoBLZ3TKotSSn+hTqwdoD0g9JUC0p4YikIkDyG2QX0s
IunHJvu3Xt1O/iFPHqyePi+cSpQpq1gKtlLTfjow0wDe+BbkLFJPxLmZ8gvDp35GgQCGlpTStUXY
Ki5WmtJOxi+I4kNLxkqTTvMa8Glyw5q4CklZ/yUR4Kqc9HWw9GbjcQHMiu5RuoGnmdVD5u7igMar
9rW6sPs4I4/35jBM3qmybU1k97MdouaBcgzRIBbz2UGPX2I2Kp7r4YmzENRdHbaRGRCcL1mstq0U
By+HptWiqlQ/G2BONpxUE5He/0tLN5PPmPSNf1xzhx0NNZ2i6tyoxSxamM1OIA/HLjvFAr+9YgTW
MIhBCq9M1m9FCZKFn5/Hdn+SGvbruRB5coJB87Uu64Fpi+X4umCLTYn3dc/6EYD6HLR7qKOMLg8q
JfX9VV7iRP/RxC3onc1ulzrIfnJ/lUXhkH95kC21t1iz0MawX0AjTK8IY/H0+VWy895oPgr4L00E
TH6FbjqWRS+8N0JZNBuCDWBuiddUsSTmzqYtjwoPpGuijf0xn0mWJFsfk4IBQMDxo7JNFoZYdJSo
cfQYqt7NGjaUN2t6m15W5ocdk5x7TeathMK63jUNptMl5B0nC40FufL4UxyR27Iy7vrU+6uZyxhl
vPMBbGCBmcQueeFjghuDxWeOUVpkYdmqfxft1wGIgZG4Qt0LQb/NGzvhu3p57jFKqVYlF0J8YZCH
n+ACMw9EoNKJ40V6n0b/agsfghER48r7lTNQFXYTKh8lHH/2vErg3Q9tcIfnwF7np3DFODfpPsvE
43QzdbVsGMenkP4rorlvO4HJbo7VqdCSgPfYkRXT9qmllOlptyHNf0Nm1yibdRxU9CguVPXE9PjZ
DWKmMvL7s74GGtzbCNk6jqLMKRU/HT912zqqtTmL0gFjwTiGpFm+akqsi289SZh0rouXZJgviPao
D8NYde8qEsAOc/vKGwVMtiUVtKAvQk2fZ5vsIaG1E0Pyr8I16hjzlWtDw3iquSiO+egR6qZmUO0J
0ICnQ9ujw+w+Fy+eGMUh3kFYsIPr3UqBln6DTs0eJBofGz60P9aQfVmf+ucw1dxn+4RmxLPhPz9f
Al5u6R3wDMuJkeX3dUKJXJeAysapAe8vwhTGNvgjh0wBRajGofsrBS27RmtL1LBevAbERC6XW6vO
+sIA287a+3DOAHKYGDLOX52urx9XvGrUyzXGipzXVUUE5I4Y3VMkPzrWpnqvQL/cVSYvHOyeqeHs
FQ6NqLN+UKiB6uiAumV9nYXM2KypzB8KiN/ODUhekEWJWHfKJFRTy1ZH/9/xwdTeHwu/FMULQbAc
6PSVXfQ5keacxzhRVwZu55dSW8NATWANGlHkHHa/Tg55mLKv5WJ7DSZIqC+e5RCN9dmZsIK+2tRj
D2yjf8k7M/YjsScyKledMGXen67ya+D0mFHTzhEAFLU/8RRwGU+wmontDxqveLGrZ4YWreHXGGc/
cyBLSrjS0qwfqOMfg9y6jPQt5vsYa+t5e1XxUaHAk/079Yd/wCPWg7hSyDMgbXnGxixjuTEOK1pV
M+/8SK5THeeQ1J0Qtk6ofTSFvb8je8XAZ7nZCfilbpW3+qui7dTpfALnfdc6Ok9lZJo7D2pZuCZJ
SKNRswPzg3RlN/9vIP+IRV0su1aSU+57wXuyOsJu+Nr6x8TJcy6YrdCefRyA4BBp/nopvt8iTJ2U
zONzGJieR+akvJ9QuXVPBnAmltgrqhsvk/9FMD/kjtRFoc0na/BS2PtqDZFFXWPk1stk/zDLfaaE
l/iH5P6IDjmkB0c9kJmwuyPytzyD+9POi5gCH34F0cQKSg57j/31Ssw9DPsTjRJ3kPMCWdH5yf/s
q2njGHuVNvKSor0hVrkI+5KABOhnICMp2POYaiUyAEqa8Sa2GBlAuAHoh7WxkWrPrjYSqNoiQbcj
1oGWOc/vAvRJOqcQhcOtzTp8XHa5OoB3rlvj49zIsFfy1DaFB0GDJsAR4mMtob4lmpFFKR9uqTx8
DPkVb9/it4ZU85M3ZZ4qriEaaG7e3E2+4IwIzmDkf7F9lojfIXe/egK9F5bGeAbYhHnbTcsPQxpe
jih+L8WWpTf5A09V6stqvMIqZC8snggiQSgnNOIUrzwaYsrulZvIxHF8FNb1O6brfz4X3C7p4HGI
qS9ojsSRPKdnDktEPf1yZDtcJ+x19R5T/rWEZq9C1GBbBLW3CWjtAKWvctLWNGl8fLAfNilLQAfY
6QJ4so65oWEJXRG4hf9mE6jOSLbBNq/pP6v3AQ8GaHU9N4PUBWyK1pNEGf+16GOnSUFDm+8Ws21H
3dA2JdA8lCUpajCRcajFAkntBCH9Wavsy9jgZsW2zKnJH85g2cO4nylGcrwuAVrKDv5NtHzPrHR5
2ATW+fXMCuCuC8N0rLuNbSFq7iUDYU+QqCxZojdk2s+G82MceAIdOrxDrzJhF3di9u95O1MmotgO
AB2ZwmU0d+RYLTYssLxOcKvpSqtxzmOAs769Rb4PXLCdnEa9krj0A/UCg+YWVcNZ6ocJFRd20U9T
0OdO6q9UUukBHD4v85YjHDyMKa/qEGpfHeAPHK8ynCyAGJvHCjWlUyT44GeOXxAMWy+ZR6du5IiR
vYqQzS9yLvWWmKU7beJNP0okAlAt7kt9CZ+kqcKa2CABJqY1Tr7NOhLSlJXE53lkzM92Llq4bJxV
5qQ6fmWWdTP8uPBHWNTG88Lsh/GrnQDJ50EVBUkqP5sFq9FNoBAjLpOqhYAWYFfKK7BsKgSfVX5n
McXte9zKKybkLa+dslvdl2QTX4FScjgI819cXx2y3UOr47GUo90FZr2I8I0XQp8Y8zrnHeP7VKXd
6RKSaE2wyMLW/tb3xDnT4/yjgD5BMODlsm4vorhmGPJ8YMaYYWS1nbGZFc/QeV+qgLHwEMmSTVus
JLun68C/1QsSVeP/YJtR1pJ7SYP4HdZOh9Yr2jNHq8O2Uo4hmSmrgwjZhgDvVt6Xb55cIftsEe1b
fQQ/zJA4JdjdT8rZrclwLR8Zz9KuNmH/tSnwn0W37inVkxMU61/hjRUTbNfkCmDK/Jy92AMbpQ+8
djcafZqebKPlEsiyI0bFATVmZNuYJjn1OuuElm99RqluLfd0Vd5osMrVz5Bnl7cArwDYtEGatxJ2
GufsKEYszeyNojiAZa4C9/h0ZLNPFsGDkW3nz8bQo5MHUN+V8be9qE4TT4o2YIadfv0mVYons0g7
I3B92bOSYP/hR2uTSmHHiYv+wuhWLBrbLGqgFP3MVZ7DsxoRgvsahaZVHt+zu4G07jX7GhqP05rd
iRSX8qZlu0w4YYhuB6jnzyprwlrw68vtgizp6JezoR3nOk5lgIvTYYadV1hXd209bx9OJ6R6N92l
DYbzEItkxV8PnR7P1Wf6GnW0H7LWzeB2f3CDZxteSf5OOQ48Gj+yazAa8MGzVlp6qW11phZoicdy
dUbDdu6R+zSQrGuHUe81ndBRPRpjhW/wq0LFI97SO3tJ0EI96ysREPmcYrtysCkoYQyeTXdUUQMD
bgEqc8bENY7h7ev8aeaKzdO4leMizZZRg7jk4PGKWPn44jJzAoWSzZLWGdiIf/LnQMy5UWx+MXRa
AhoGBkTAtON/yz2QLVjo70l9GW5YUKG8Mj1/4Tt2Z9YF94T4tZhpwp6ce/IUdvlpzZDVqKh2RT/I
vJnZ5ML6XE7WClN5khFBXbtI7DqJNO8LP4LXe6d/Pls0JlWao+9enQtggByAyK8LOZyYwWkSjSFP
Og2ii8yaOb4B9cOUTr133kup3UhRGoA6u24QfPENv3JOp5n0VtsKbr+RVySXuHwrVSQ7mJO4yny9
HBDIbpN05TJt82eTQ3As18VO34U7gxRavr1gb9rdigxXsq+9HfgVGOYqBWsHeUb4HoPpQjQizYYx
aGGf30BusbDV9vuI09mTLBUNqowuP1PYEVAPrdXOKW18RM7VGRt9oED6qQpWRSVxD+ngt2iVGAXR
/K3v/dD/tGz+WzAafNQ6jZRn+87SgEnnWMNAAN6YCLqJAh7erpUDGOahBdmqTQDa4ADDI+08B5Ku
mcC8axF9o4FaOqw08fGDabjnpGf3SwHVfo+6+NmR8h93pQCv798bVCbbx7YTcHkFydHrNVeVkka7
xgFEc+fN6aUTvfv+Bt1H63TmnjlLHU70o18s9zM37ZtJzRV1eCv3id9rvh0mFwFDMm9YjaN7Lx2s
9RllKKIt7lEmYKYwu67PoSvlIdfWbbx6au3xBNaQ5R3g6tuiIrRYCKFAgTpFW449QV7ZHffOFcXg
qVFRoYO6FM0c/9OIBjI/vmMEE+2daxH6+7qVsouA0oIgzB/gGr+52cGKQZ45gRLQTyHkWm4iup3N
/Eocss61HdoD8Zj5bXOI1neuc2YvusMJF/ecj68Pl2EwPekUwWpTrAQTJsOSOb5YHHTjFw5x3QxT
GVQnqrFRDt8i9SjytgZrpoyXExfqHac2k+KW1VMimj/F6EPiKBp583vQ9JjeBeBd1jlSOd3s6Gqc
fbJutOqRJUjP8/vjPZo5AHNDVaMXjf5SENC8iUpl+MWOVcZe1bcqQW6JZT7I1ZBbq6wLJxwp3PXB
QmDrPqWtuBJ2FjjVC1mLbDpm+8XAx+5N7H0r/4AgovGTKZpxkeAEYDsRPA2sddFpAzZk1y2J7Mfq
UJ7cn5GscG/Jj/WjEaXtn0tVtg1kxV0EOevXzeslWkUCGwfPx7RHEGiQo0E4U4l4Vaml9vqkGeaL
J84bThOxEwerrLDuRfhk/imXGB/weWkNggd3B7SvOd5D73K9Ab2TvkvsYpbYBtPd5D1o+RzdJqN1
emhW3tVPeIrkuBx+9kkefCV4SYF2vqqs7r4s3WAjN5Fo5WvddKTs+Ap6czSms4alsyz72OHg9RGv
dSsB0XsRPUwOjfSXIKNvsnJ447ZMc+T4b+PbVHDtLZPp2tG4xUMFT7r3pF/xeeBncehMoPKcRwBY
zHAysPpHobjRFoOTWGlVeQ5VQzVxf35phorGf1D9BEdTnCK0395JFVsKDi3rzf35BrLapeodKSIX
b/ThzAQ91ZnW5G7hkhKEjIUbewZWGntG7XsfXkL6MtNzeVUfh8GEzDtd51csUzG4CFIUnVk5h16+
+guOVA1xe2YQjoHKmkCAYxqP1AumolT4Ezs+MzD5yu/y8yi0qkJhqfRUGiwjcOUsxOQiEaAzoXba
s14k9sDWjXfY38MXzQFKDrIl0hgG26I/u26BRlIHrnI7nShwE+6Y8btSbDo4mYfJaE21C43VDKTd
o7CbJPeHCO2QwkLPDYe0/GQJvnXvxdapf4dwX1QuacfpIi6Uo6umZWlVOYJN6H6Ef7skmXuIRoHT
2QUkTfLgpZlyvWbp9xdetdPxz7vxVNOfTqNUsKhqIi9kzNAPOAXiOKnSlmpIrCkcVeKEs7zakyQf
WR1rfmNC+Jo+nAU+jfM/PfliUhRGmuMw6s8VicHprP6HVswTPj68xEzASPMgDrP0Xuau6W9LMr7W
Hak7DMBeTlaPK0bvEcHU7qWfLRxEr+UsuLGs56XfRYBSHyyfkWrQk2nGmmdH/7GST5mRQK+EUcWF
soFRntpZsXzcV8bfaTSLxI2de16ffEB3z9hd5F6yn1qElU6X7OiJ1x7QzLmZCrcOE/R8q3mO+Mqt
ywtM0f3U7GRig1VnoVFdoFexaaiSedBwv9IzQ1pIwqWntyE+YIGxtve0GXrrv8sIgknkYS5jE5DU
b3bhOuo4csDkHNc3OLtcgrEERyT/rv7tOPidhr9+wPj9TJ5IyKHurSypLI/MAzaXShxkWjGwgtKe
iYmVHplhexBto8EmTSf/1Jznr8vmoU50EP8EvFSVIjZkuB8QcmbP0kn1thHJ/GUbBUByqRD+fHG5
1IGNoD6b+8Ygut+GPMb3Zj9vjPT/ZMasecKngDCyjG1CP5c5QxxhUH/CdvAh9gfxdhmq2v6B+yhB
soKlh2NcYgge3W0YEWzxMiVa37bCEtvkALwwPqUoeUFlVlNttvSax9DS55tPd1m4l7pcRMw4mBPm
B47VmhLql9IMCDLolZRyqCd99ll5ghRPmCsaq/zxHlveTKJftEN4+fKjCMPjiZzfv5xTbHCdEnlm
g7oZZmg4jNKXm9jAt809iIOujJ2+saEuZJYtsnPcq7utcxJhR2O0CvRs6QyW82tTbSs4pvB99w/t
AOnqaWeCQoCXuW+RUjMkI+xp5cTWAhYllMWkFYYWz571xm+LVPbIY4sM+t5AwWszYIXlQvdD7KwB
b3Ux1grxVL8gSoBvEH20I1P4VBNVsJNlEKpu8iKCwRSsmy1vssS77yXebC9cVCuHKsJcCFwYlycU
1dc5NoG7khu5/01XqQYewRBoGH1poVSqrEyxsXEECa6udOe/ftc5aQfmM4+d5XuR5fJbb3dx3Wl/
8Hhyg3hECn0s8eYAEUKfDrAXbXZcZFJN1xYiY83/xk/eZBK6sKSHXxxLCM5TmBOV9FwMQDPrwM9Y
Z2d4In1zX2Cq78pBBKeo3n2sFhLxUYWL5Oox4+ZJq7JLGiMJI83AJQ4ZpYHPWsPuXsuqPnvza0pg
+AAZkSe5IR8pa1mDxiQy+LqT/Nlg6LUfguAKWt4e5StqUQkFNkf0SoiGr9oUhDIN6g/J89yBc6om
+TJsdZbsZX4w4tRfGlboSq+9PcIUmgwfl/8vFmw5IusgNtqIhX3iOtlpzODJc/DQyILszZ1srDvV
77KYaqARcW2szy36m9TxMOZMsXGaNneiXV9yS31xilLwO9xV62DmU2O2sX4uCWW4z8Kz/lPz8wXT
EkXsrBoaiGEaLPSz2VfKAdiOpXoqBI63PdBXpZZe3/hV+98uv34DVv6S27aRZ1ao7y0VNq8UYLde
nCnEMIU2BedButyYATxX9h/QQX1bGkOuVnEGKNYUFe9ISvCSJdiI29e5cqi9orzKPLlxk2kdu0LE
wv8WQmUm03Fnbrzh882OQdz1P6hSqCLoiy/7WIic9Ecg0j2Lyvl9IapyAVfXltXuRnm9LDm0h4WZ
KdTKonOWYmVHaTpgq9CDX63Bqv/EqYoI6BsKgFUKbBZRq5ewMImymDJjr9ylSUH+iJat1pt/pBx9
WXBm3pB/V0qHqH2pEr9ClOMjiAG+SBjiZiVBUUz4vaD6PMAv79992smJX5GpHlZev3skhsXVqn0K
ZrMMfzCyk3vNv70SgH3fnEPKFz1Y+DwLGhxLKP+/GlkJzoPYaOCNa8RrYbbq3LkcibOtPjeniBKS
CSRIjg45QfEyMm9eAtPAI/8O2miApO/jp4Q9QFDS6xsL8Wrdm3/hG+BjjMcIl9pdrXGtzd9xsmn7
FBtXgClGGmyP5vYzdCs/lCurJ++e+s/HYsH5yanNZcboOgH9RP1ehGBx21CNv+az9NwsjA7tSOAm
KyTcUM+AH/yhQuYIVEtSLJASOe3xL+aJlXv/xkQMwh6/9Fjq/53MUEGf2u5a4ikkmnBUMoJ/Rl7H
88Hl4QYAIkLbxu9ux0Z+LPJ/8vviyDp767tMLxstCr3OgtalQTGvGyxKLA1tfUF2/HVpz96fR0pC
1uAxFHHIJK9DwHw/7JCd7bxONXGZ5e5Vm1hgdCJFU4PoSknWqgoJvppHYvq0jFla5LAdRvicGCZX
fMgkx+mbZwtxYAy5d0vyht3yNf8vGXFiTZiP2xhqdPcBi6+q42OwNEME74rONKMdWAhSTY1+RRDD
bATTSVmxxA9ZSb/53GZbw1Pk4Rt1rc19UZuhY3FNmZQHNtWKHtxR6Ernt/fnDeLKOIl9NE4JapnO
zxS+Q3kDMhMKoEtqvV2HCj5X8T/PKUASP/js07VbFt6+4bCYCIE71QMfb/lx+bCsYjmatFO7ull7
4uogf/X5pUK37AxY9iajyGpd6ZGHdYAd3v125R1RmOZlMIQ7qsFiIbAu6fYS7Ro+Vg9o4lceiUaU
9y2/2qqjY7qUBk8vCHUiGLGRBEBKeRIzkZKhXkl39oHAj8oDcAB96yod7KYrcH9SR7GE7MA7iAV9
e/S+90uc5RohVeu9Yms23qUT8amqjIh272JNoZx+YlfKkXn/2SISg/8Zj+SOq5PssHZmB/wNzbIz
Ob//GD6z04lPqIo84sY6cs/wX5lDL4vSwVSxoZGRF4Rnmx2NXnUYWTslzcGhsQRFAL+Ka6VhYneI
Dy+cHEvLW5ovgq0bB4YaT58keLgdh9Q0rwXL56XhAEPCVaWFO1j5vHjcSB/gDOqEiG3CcJIfRJl5
Q+SnN/O+pDFRZvv8zR3SXge+EV1zItE0ERbl15k8BoqGv5VazT9PKRZyvtWCebqsxuBX/szd0bEE
zJwmoBdJK5IL48KRvL1L1LuJiqfbl7o30qpgsO6cKa6/2ycnNRqzUDw6DiqDOwlceAjQILCTs6bF
ZfQWof6MPLdtzf+Lov+hKOAVQ4JIRm3QjMs+cAMHPmOBDDmHEgEQvFc5Z7OPDPhlPbtV2C2d9FA9
iwoGKrTS2t39lYNe/ASnIIqHmiKQg4hvpjNf6ERLQ3aouQH9ng0YTBeJRNJsfFGPLtfOKZ5pHUR4
zRVOM9wHyL3RDVgKxlRcQuffB0/izXj6DkR4YnGSip0IUbGWHVsLAZg34+uT4i28h7Z63aoOYJD0
OpUmL1FkMxQGoGippf6ltmrmXx3FMXHYx7yV4IDggFir6rhav1FiNYTqniFnsYtcPB8u4ZSJ59Is
Ka5XKG+Yo9BuF1/wu/iW/g+boGsV+q57YvP3ITYJjVr2RmRRuwLJG+0DSa3yWktPnJDB/CFyQCss
UKrRv5PwKqpwKBSuxSv0onrflwEE7saBlq2IbSANMEq5WZIL5dYANkqxyIo7teQEEWokw25HU3/G
xYwZ8CPIadDIWAyWWQxoVGeCYdIkt3Y6pG4FGvt1+mZm0JB7Mo6f3c1BpirZOY1qN1YjJpedDhpc
kbgP9DQnZqWT7uNQHwqddKwcIQL23PIHtCNoiSmUFzpwmBsVx87DT7nDGgCWhbWqLgROYxq1rvFS
aHyq9K3JKQy59nPbDHgSqmiWpkGafQc6+qWXZxDGZLLmBUJ5X1dun+yPokJs/vNOKhXnxc9Hioso
i+coFdkHz2IVaPMcSQmQzhr8oKZmracvd/4XRryQzFyrLtwwS7SF2dba1cQNS6XIQjROEzjK4rY4
zt72wdDMjdN5D4udVo0ySfovFYB+FdBrXBB8OEQaUnzshGeOUp53wBdmhmcuokvlz0KuqX+KJZvn
ojjpE0hDN3nZn+MGX51yE1/dHu6LDbqflLDmXArNl/h3X5ZNFyqKzdJqK0/v7np+Ou8m08VLeJgW
iIKzpgQuwRek8//hMiwohf0QHqK5nXdovCW8qdq24ECmj0H0nTzAwrW2Hx0UklJ4NwkPtU3gO521
Nt99Uf4EQmJAcUZ8vqlbGi7zNRvNYpgl6UxpwufuVEqgTCKbMIiYJqTGuZQo8OjIrQhoCJV527RO
fNVlF3pvoaUm/rsRZNXuvLdGJHp4ZIf0OloJGaLaOc5DqW2AzJgyE9FHRsmLlznBWkwcpLLsB07r
GvQuAzKma2SbD/G4HwmCv9U9vxCglU2y0UAKfuA836X7NLAPrA2SlBrr5k4qwhh1ZuJLuFt+LvI6
tb42RNYbohskM28ID1eoRMibG7VAbX/kjcx/gpZBezkcyCnAd0l0jOhY0x5mVyl/V+7MXRWhgGjG
7NfI/gSa6Y0R65sj11dWBudHkH+nMJID/4V5QZOb1HrQZbKiOEMKVwf5tS87HzawWG5HSg9cu0n2
/M89+/7o1G83prlkhapAKzRF3WtdPJtMKCNOYGEAQ2KHsQmyrOatRBUkizvcGmKtx83s8CL2y93B
DJSgjJzpQdB0Vx/d5qD3cwhXhMiGEASGHMlqtZmYExmXJhInXq2vsLuA1vGsaDmiW+bX3Ker0vWE
qZ47X6Pe8vPrN3VWSm+ttw6pLLr1aJau092Sln6lieUtjTHcYKcarjpLkPKqWDABIKbzM+nht0f1
PaN3/seJfuURIScRx0OE3HDb+4Yr91p+TaXG2lsXmH3bTX9zAb8/AWQ6OhlQCySoJlVGrURDB2Gp
HvibnFnZ6pSU1g8wE0Kd9agYgvbD5zGRA4X9D49ulav+hCQVQE7D58kkH6WEQdiXqzu4VxM38LNo
z2cwbaOFy/MK2sw7THvkt4CVyxMPi1KuYTeSKyveDN7E1J3iq8lYrGXExeNq9KOf2nS2yHRhmYd1
esHd4S6VN5lYq5o92I3Djac5W5nkiQ7wS/1V230SDycbgG920lJ2KzpvgH0bl64DvcsjX++CQxUK
6U1SMFgxLZFnvf1o0fz/NXEuo4/6HqNxGpP/OF8AgKK9zVUrz8NhRQWQWJdy8SUpl4Y/KScNU09J
Tuna+Gs9f+tCtifR2Z646PhWo6n412U8+UdCD/3EqMZRIqrg3CaXCHpz+3F8utH1OkjB4dW9BbiQ
IgiNRx53b5GzsGBaKhtxBtWLixHf3zsZEFyijbiKQJER/LR7H8bX7GBjjE1JO0yZurhUrtakGUdG
Fu79jRTXEDZtPbQ22JniaEHoJg1PytDZDK3SmUQDiwg9Vc44rZLGL1rGb61DYmbNd61WDjFLzbfn
euodA9fwDj56lxt0WGE7Hzv75V7SlChi+KDVT+B1/ksewg97fue+4nOa/uXrlhi/LTlK8R0Odfzb
qSPR2OkED0c2ejmc2QcLoABtblka4UizKGR/aHdpEyvlUh0Pd5LZ03vTjmuaGgqzzyCLg8h4HTnY
Bf125A3acbFk+4OMPz6K8mKfI7PdouUmQL1RikgLmh19UzAZxpvaYponACf1sCriP6Bc7702bA92
pmLLWbI6Aks+mQQWsfkoS+Ni0quDiaKYoABz/wj3I0A/mv654E+kM3GXm1BPW1YP/h2zDh5iVkhI
FyzltS75xQU0FylbOmsBlxlZSdcp7oZeEyctmXSwNgh+/6sUTjt/zWZEhQVYQkg/3G/wpfmGHf8m
H/UVha3KKI1CBIQLru5synlIGUTlq6h8QSqCwF5Yo55VKukyZ6wlW0IyYruEZ2k1/wVvmOt4jcu+
l8k1XJfpWinAPSSbvLT7rYC3/gNCUC8LNG62fLm8f3kVHtNCExY3Yea7ZQVpX2Q5Bha7jEnLbPBs
LinVbhsYrU3ZjHY2WCASCuZN5H0HlG9zbTR4LIdhY0bE1OcgdyAhjw5kfgYj2GcbBCugMDLrdNZ2
XuTv424l4gcyhjaYdSBOPtT+4/k0pUpHV+DUJf4p5inLDCOyrr5qiUCjHGfSAgelscFZTea0yIvl
HUNVkHuSEbI+w4fo/6GK7AMe9rAW1/jlZrgaGg+6SL2xYu0T8jZbbypKmNok1I9Qz3Ax97fvXjrs
nWyKEWNQCFqIAUM+FCi/adLYHFQX0o96n7828N15p5Fs3HYmy+OEJhw0B0gvpjtUA8GbRJuU0IO+
5EjaezTCZ7AVMl2kIM9SoW90Q4F9i1/fETgtvzOHAFmnjinsLlmt10Si/15LJ/z39LE1EmVT8Tjn
bReqlbcj2wYfM83EkBnmStLcDaARmKtFjo/F+8BGD06E08RDjfpSgL5cIOJUP+gbd9aM4u8IQJwb
LzqEnDVpVNEPaRUHw1kGevVvVn3BD6hS8XIBKl6eh3LsKKDPdE2YM4BHWEW0qbEbq6k273vwzv/E
9E1nKr65w9vhh9/Z6AOOo+EeUlKrFlHjBcvNRk+o675AyP72h3V21UmSoO7lf3CrjAZJcTPdM8ZE
V5zrkHa2uqYWc9snDvN7lIca7xxXveqKn42V7QzMZ2j73XKPXUKLfK53jr6OF5FyiVvM23RfnH1K
OhKiJGReKPanebfhABedtZhWnxAcTejNBJZgkywONTmQ0ATFmObtGpyZLDTvbwrmsOvFfSEhHory
aftjoPtJ3TcE5hQSzbwmVkAcLUl/Prxk2iAmsp9vnwdV4qa1sdK9KiFG9pML6T12MjVkKDvELORv
MQ8uiML4GJGVARCrKTQWC7WuOlqXeAN1d8hhFdewomQwdNiFPgVxrnMII44+XyGrfst17PtxwLKR
HrRQrMcspLy6VpZbDrw4I0Can5u1JfyIQb0AyA+bkGS/J71GGiL/GNFbj+eGUdGAR9Ypo7q83SLw
6HgoLi3rzRT2A/fGXXT/J8XNlLlrSMR7uZU9ydbsyawPrErYGSuNacsReblxUBZfp/sCEYa5UsxT
tV2lVyNy0FfnEgpUhbI99/4bt8IZZRWc712z5mhNCN1EJGamb3UehP62zTJ07mRTNBX/VYcvk6mW
6GWb2/yeCQPcO89QtJSy0mEBLexiJAWednz4lNJmURsdpWzyLY3j1YJzCQB7jv3t3eMBvVfcnjrW
nT3moaNPGrpFLDWSdt55liLevjLhhO0eKBiDoRzTLPPFklVvfAtKLq/Vx5grjGAr5dEOaQYmnUUM
bjSQHjRpnOrhFwTIqgGDEnI03amNn/WjyMGIpgV/qmq7aGn6hjCEQVkwgHl6jMgYR0hSzTJ8nmq+
WxzjdqTOafNrrKLtYOvIGYaE8vjgei4uu/LIhrzYzapRBsg8VSeZ4UUVI6D9uaovEeEmJzbNx5SQ
R0tWGasS2dmzmhxyoC7tZFMCjzYPiUNnXIZFloTFyJa2P8hV6YVRQkOzt3T3r1vhO6sahTVpes3w
3aucpp/YEhNsSrUuhjOOSyWB3oZ9K2ZjcIMJf0LCmM6ZDzLc55EBHXQTHdumHEP3K14FlG/ybBrR
xgVnPHRO758bQB+DiK2pmt0cXzEmzb/xFw0Pyrup7xCOUfrqPMoYl3QSMCfs8fqyKstOf2K79ofJ
JsRRnZQxdgXmN4kx906WJjkAypAv/itfDWxQfdRNPTS43v8HiQOjy3l21V8DaYiqcWeP6yvo0ObV
17bxI1U0r1lyVo6/4/6SFbXPGXIGPLYl+nFXD048gF+srmFUH3GohLntee3og9W2mrHhGQTTHYKz
+ldlaVE5xN20Q8JltrAqt8WXPOnH0A7xMO+mhzVaQ/85zk4RROkskMoRPkM1HRvo/0m/jXE/FJYs
kBPmu1+ZOyuWe8QoKbIi5SYsU6l2enQEMptxnOVIo0olPI1Ly/qYxUifB+o6jcrettlsp8e+jjgK
MbSZ5Tc8ihdBlFLUs8loDZ9vluhWqOrWkOefz6zYG7QNN4RtLUY0T+yZVyMFe8M4USYgC4v8OT07
AoKeyr1Z/x+hpKAzFRZANMB+KVoGsLTEnWfeFb+PEZp6pbO+dQ88bJ/z4dHeQWDXL4m37Ckva6Ty
6aGEc2ywdWyA7X6dbu3Go8VhTOguHzzo+o2rrXg9Emj2uBhupYaOp46cCrZVTMPVDYVOiMgblXCz
M7VWKqwpHJV6uO604iT3vNLcb430xdR1jmVRDUJchurbiRFMLvUvuqcbJs1DXveqWEWeU3wR8Qaz
+nKi3zCUhMhKI8TRMr/z3iWSIXJHYM0wQ2Bt3DOl3AZn/Bn7GwswC95L6NZvfTmfXuhXSfnVO0Av
rZwYzknodyJQ+JpOlvFCofhnF+mBXMNdsvMl0Tl7ViAQSYTjMrm1oDxGZpUbixWStY1ZL20t2h/G
n0OL9jS0vjLgaQ8SaAqvk+hR+6VICdrI7c9csX+Xrb+E111m1NjC7mahxy8I4I8/o+AmyQcF4+HU
7tZVh33+Muvigm22OGc/RZ2S55MN4KnGCouaUiW0zI7WA0ixfJFEOhn6r6g9ULlPIdwEYgGESKQM
RVCskCFkxK3Yj4V5ObYyAW4Oxwub0OkH4g/cxiJLo2g+g3vXEtXfumkhz8Ck1mEDTVEJrR3KVXxi
lR6hlfYPPSRsE5NYRlrsKfiU56X+Yk2guv26J8qJAfTSqxB5sCNEhHkSuutFMYFJwEJIGW5Xv4+O
evIxZoADgUC1RRS92PNASC4dLXczx5ERgAknXF3GB4OIJaKCbSNWrajn6rJb1pqhh6lTbc75JrNu
gUPTtWB4kTIdEOpo79FVl22nN0ppQ5FZC4zua0uOrqU7eTl8t9WVrHmqPoN30YpfwvkMFL3Nhsg7
w4MYQ11X0H8yCG75Yi30IrHonO3nQGDnabVwWAmH7zVcvT7itMlxf/+ek9kNmu4QqZV6/nDYyQn6
MPlwh2RyfLEIuCCx+Vfidvu0oGn6F6EcN7k6NwYxN2UyszD8Nk2sE2aCED/LMbTdmHstyd4m0BCb
xfhQzit/kwAqlBy7BD+cgu5plaaWJmHqz+axvHF2FBdL5h3hguNCf8Oo3NZsk9oXENJh1DyY4ca+
wWwUu1DrWpOh+HutY5lZf7/z4biRA+dD6TDr3WOTVhE+p82lFdE87oWciIlEUjH5iO9XaBszq8hq
o8Y4aIRqUPC93YQaLpUxIFHlBz2TwE5HaQ1bX4D2MNr3plcr5CXDKwU5B2c8lKn/6p0qEpVSjct+
juuV0lknSDIFWeOy6hqUaxdLbNL+aBIH8Rf9epTEBsnM6BLQRj7BZwhl4CMvjTUpWMwIP0jdAFUB
g/7uJ9hfLe7/Of8jMIUfnEkwXTYWSf9HH/CfsNsHuyTpToxUT4rQN+shrQOUL9qqKt7Y6Nr8C6Tf
oGUkroE2CmOQgwMiRhskO/o1ONN+J5+bKWzP0sHOHlUVOCfpIqnyuWx/h0BVslyBGAz/7M9TsYtw
POiwFh16P5JTyNeUrIiLsX9MKxqO1KMv/PLn7t4etl40RFrIVgGFjl8h+xbcDbUNFxEeJsKe7njX
pTGWivgJHkbzRMK4h6MvOdf16paiZhvD0P5JTsTt+qqsmmIK8WMPUJ7yzese5Lh/3JQROOD4mc40
hFLc+R2FK7a0QzBGXY8YDi42kPF4DhZq8y2mQ915Xb6N4ONlNybaVW/Yf/9u6wEOTvktRKveZqOI
rR+SVGxUk+XZ6WHMPkr8fWaR+3pRH7zMm3d4E/Vlr1EYZNEEF7nw3IrJzhXFGh3Bd3OaIQCC1ski
dCt2Kh05tEHG3doqOdtQdojmTJg1oYjbhkSq3aQVi2Fmk1i/Mm+vV7BL4cGkxOBT8EBKJVwy2q0y
L69kuVIGbSLW2z9rVwZnc7VG54z47msO1XJdt/gutqiR8BE6eXmRp75CagWS1aZ1CFhJnujnAAQx
/fbUKRqPwKaENA9b/5v9oXODFYZJmqP0w3vyY41hlkcGl8013GAO3syRAoP/7aYCXlcToEivSxrV
izejvetJR0oyfFO9tPni2itYnu30zqaqYWmq8PWtzzuzNQTwVdp1NE+AGL4A8HomVOKgWgzdQVdh
iVgF/lnkNfUzDlRCNF8CdFjc+ysIRrFJEjYNKPzyQ+TgmHVFG3SGryIkTsx0PIOSs6IzbjIpaeVf
YH/Cf56Nb0/Zk6Zuha9C0Gc4iUayYyZvitI6uBa2uaoIsQE9yUH1nYuxuc1rywu7VwauUKAC/OM3
vK83xbFs+3Pau1JCilmg9fsg61OSiC65dvvThnR/rWhqrXeS86FR8kw1NC1xXA/MpQwrPaxXrPq7
JiJEqiIRzsDSpK1CY974jWkvC8J7kVEa57wrBSYVMwfo7mTEq5YunQrmJPDDtEEH/eDE3RPQIlZv
KidtC5AruEDUthkIFb8zqXEZtP4RuIVocu4lnT9A6eQC5Wmik3kAlLG8lDEFqZ3qE7044IpL5XhT
WvXAd/2JiXd8pTlR/5HWZHP+pn1VvR9XsTTUhzDEpCzqfMHv2OocUk1ppKHN8P5iVZ2E73XizZxj
c49UASAnCqFhlfBABb6tMQPevOPTvzjnULn7L70X8DfngDR2u76pkCM38HXV3KbCgAwzsmjHOISF
zr2wC8iXQE3IKUTZVabcrd/2iOS9XTA2byG0f36Bl3G9rpY9viw5N1zAL0syywMXyDHY9DfFQRd9
FLiHYAGHguLe4QC8dEpLewj0BgJWS2ilKNzy8EHAHo0aqdecLDVqNuzUnHw8cC3VETKORJI1LzTw
s+l9FSA1C0EpTez56ePejY3ov8Zy8tjVH+nT79Ugqjqp2g1wder9jDdiJJcHmNmq6NKCAJJISD2L
bRm5OMNzpEiw3X7xFuzGY+pTIRlSyiGsfHG17x0yoMaCUi6Ria5vqMeaf9KIztngij8SX7YB12MK
9UDg5HMVa3MhCfgs12mRdebyLNATmXLqhcyuziLTWIxZoEGsebsRKRZTiCBr+CWuB/zEKddgkmdh
QKF2xjM/Ev9NjAiEHtG87VKPkBl4+11HkdV+ILUbevIE2dccTEFNfTnv/KLQJzrYDYHzDfPuSqNh
va8qRb9hyphHyuZdGaIBYMZiFbWapUFBSfSAoyupAXlMeWWSToPKKiRZo3Y3uBypauvTKmDyFdCg
R1V7l4g4qgl4GyLYIEZgsLSegnsAf2Os0OPg+gyGPLrSFTbZWb+X4yLfRm3lD5GbqKDZWrHWRZD3
Gmgu6d85vCQpX9Y2LPtbz9YOVbPO2Sx+bQxioDEnuPRAG1K9kpJ4OFH7I68xqADo+qvqgoeojTZK
PYMnE9ozIzL7eH19J3544/3Y591gp4T6AHDVJ5ifrNd0+5QiR3oR7MzvuJ6IEnNxFocTJ8QDDzsc
h1kL2rhULK6/0T2LhjxCsfZ3/FetrZxI1oLzi1nyfcphOvP/HcdZMlr+PplpLh2eG3iScjzbtqDD
tqHacfUqIAEtNEXxmN+Uwp6/b7oj2xA2xxSEWq33LAxlrzKTe4l9Eom20CMZlxlLfRaJQ1Rw4X+z
mHiMAllcWojvi9KaQoFXkv8JY19AzA7/kJN2sLadxg0fc4O8G1e6Y5EcnHN6NcQxzH35A1epkjgG
mVz6miLBO1zlwzoluA47/uy+FBp0M1bm2P6Vk16wg3c7Uhwnn6sCC0Daal7DhLSjWiQh6yHgyM4X
7SMWF5CVZ0q7IYT2Ph3EYC7n8dqzDUW0FJuep8MgOB7/WxoaQnUgRxUjPd5Xrzl7o2vuO3vAkhFn
qMRd0y7sVsX5d5ZSo0ChUn6EmFLSPaFOckWUEcKNtgINTS8E1v7RTR+5+jlhW56QXjFLsdl/ZHCF
EOWyNBZFzkfnz1t4+/XZiWP99XuUoZvFATwNrU2ItZKLGBd630d+g8JxdUBNVv56dN+ohz3IX7uI
xZGASmFshBN0cILG5bwEu+vR9c8zhtndCmsp9GW7qUr0LOPL2TQC1uWid8i69UuShOeBdnbLc3AE
Hh9iyfjXlZOe22yzhwHikRYrHUA/Yw1tDPiRLkPa5wZWbW6XwgXIezh/bu6waJl8bWvT/qxKqItB
s0H7ibI9+isQVCI+uEeCOIugXHSFCaxb2ytZ6id5Ud4Ji8TXoi5hgS5wM9oD11zUt8f8wnvkdHvW
ILVX6OiDlr6BPab/LBtXJpvPBGxbmeHrPTBwpnBLP8gvRmR5634LvDUnJ/AanzKWKfIdheyngXYR
bBeWoLolNZ05aWiGC4/8krqI+oNkdH07B6K7sKBNTLvJZFa7JkSOlBFGd951vIskxQqY28PT+Z56
n/u23YZIOZnjyolYb4ypB/k3N4Bv4ZVSbUPkzrz29HSprwK0BnkQmy4e5abDKiui9l3BckqN08RQ
MOO6vRsDvgijS2cM1wv4uF5tVoVe2senOHikLF3nO9nOT1bnLyhuYnBJPTcSOkqvhw0EPHyzbaqN
og/YbAEq0slkdF7Fs8vOj71ZhEgptm5QUUFG3ngo6CsSiVh+jjKInhzNq6nwgV3FSg1oasmE6Nna
+geugqB2Jaz3UmVfOFdK5tzBmDsYPNsy391hAMpdzqhSFSUj0dsZC/SQFZ4cPfSkKdHrmEVXh90B
K9HHtqaMW/oWXm1jonEBbw54TRAVdm9N1AxZCSNiDdxWcQ4RoPvgdCxm4ZWsl/pHmcEvQt6CxVO9
kNDMZGaIO1e89mDA/RkK5nozhFIgD8+nai4wlQOG7z4E0o0/74ugW2GpFmx96R7td0lHJoOWwBcC
iBzZYs0ZK6hOhwvwx/oq5awNN6dZADtI4EqeAr9j3usr0nX8Fe2y9cY5JSdOhNSHGVUVjmrp5m7T
QVMLCkvcbG4gwQD34+jDQcbisgd7JyO3Ut9Qn0AB/6o8Ksfx5i5QdHa0bdXR7sw5sSxQ1AaKUnML
N59hghTsn6ZlXCxoYrdWlget7I72VRoNJEvcrfnT9/gT8LyLlulQYeybQriV2GZagNnEHYxEfzpe
sBpDwIcmRTni6R+RmPbptjVmuOHyXG99JWpg7PG6Zkd9RKrTCfXVIZesZqnyptaroMxMOIhq9CB5
dekeHBW5l8IJP3EraM/zYQA/vmOy7kDp9ZBIrDUJPdx3D9I3fOOLkfnbpuBlTLhbQebjT9tY3e6h
Mgeao/lfXERgAcB8GTnoxQ7kKFSCrgETp614db4DLBiL404i8z19Y3x45fB1iyv4fMctMf88JME9
p9wYE9CmhTzzmyo3LXoEuoHkbuzNVUTP9eNgScvFCvSS8VFj4GCMyz6arVVOqLnLRq9R/k4oI13W
bQu0hx3EkLleenGVmD+YbMGhXlJ3cWh+6Qcye59LgKnngYobyukMvGYlqMEcd8tRW2HF87Zsyotd
XnwdT1zwD0ZFKrheHAgA+QvLXvRJW5ENtYMlNSGb6g7ZD0iL/Rr7yog3OQOhfylk4MnZYIc7gtsp
2lH570Td8P8PQsZ8rOS/9ZSxHPlzmjb9g1do39WmrbO726fMYT6/VqLmJRgPaCJFwcnSumgzlI0A
qNunda4BnYb25Eo9QXf7EAWe5i/bN2SfEw3LtHuhso21olSFdmIdcUpOxx4s+k8EoPUSXFCwJ0++
W6zZdVEhOS+46loTD1VG/c9SJ57BjsXlIPfUscPG8eN3qNB93yYb68ENQ4vfvKqj8s/CVbHXwkMp
BWjpCk69I6YJyG8RVtZeTe6VvKcXVYvlasPYkVfRTETA/pPC/CAQ5GxQ+XJgc1s05c/PO37zi1qQ
nwrHIx/+vn12WjpqOjBlWzdwvr1sP6OeCHeL20lMWSHFa/h8emG4fy/MZLOEmMH6MSYQDbtJevWj
ZHgwON4jX3KeIb/kwNArBVK3ca5UGXlw2GUAQC+w4qF1qLXrr71Bz5NmHIbMtxYGUrLCK9WPHs2M
ODqZreLK/96bKVaAoCLpt5zdETUwNFZKTF/Puu6/ZDmn8CZcQVMOoAhvcj3ItuFkN3KRgkumEpfM
Oh9khdyUtoA6TvJNxj+WRBbi0rRtqe/YQQXpwihLaflfJ2z5/9KCxQ1lwjk3+hcVbXx2QKrzAeT9
SLUNXaydzCOSJIq2MHNUyox5thHYGolecb2fZb4BukVN9JBpfDjwcR1r75n+uE23yJO6z1pjeGOS
TTH0OyItB1xHNc6M8hWZCh5wvwYqO1vEHXN+QYEDpbAAeWa4yUgrbNZ1S5FQx0AXtg0+RWe/8CXo
/8CTspYDT6Hw4EvmProOl9qX15ZrfVj8fDQsGeaqYZgMzvSyWDsnsgNO5qKxbmohg4dxXV1/Dwcl
qkZpoj5sPhB8cKLmnaTNLNp5Hgj0Abu5+ki8S/6dHyIkJMxpHgtqwV8wjT2cKOxVWhiy2bCY/d7K
zF4oON4g4i8sle62mrAGYN1A/Tqa+SFlFS1D6SwAczXhF8t6jEqVd5ddMHF9vUsx/OKaK3wYjqXM
Z/I6cwdpk+Ch7iq9lcJMlzr+VRQEBfhnjOG7UctZ2eZUcZnWriLKvdu7W7UcHZkctgratRNYzzOo
2YK5FUP997tF7nUl2uiJ1QYxJJAQ50+LIwFLFcYjq8qjGBQSmzx7isI0Ks8fp4PC9Kii6g+ggCG+
V2hn3n0mM/DZ6yRUVf20yEAgJL6BMrzw9LvMsacx62IGp76MRnx1T7xIjUQvX4fSJWno0niERVH2
2miaVAumO7SdZ4Yxb52Y5domb/ZBEvm/FPSwdYXv0RjTY0lsLNlFRgim0qi/C/SS66eckUKreYXe
euzgV7/bh3Mu4b5/UIXmcbl+ULsOQWtDGKsvzRy3Psm2LanVPwi0ap6H+qwEUWsd/x5sZNA3I+ph
H4Ltp7jRKKHZIxoIfAijnQEzbrx43ZeOVvYjTPeiSCeZMWlIj2XlzdEkUn0A0jpvNSc6e4RjI7a7
R+RR4nwhFv4eaTtJRBi+dnYqMBHh5TrWrNKHnbPkBx/yeI2nwXWTvPsSo2mZ2PxBB/4QNNvKd91d
YDT4T8xsaIjPaFDq7koxiLHrvPorni45+PndFUDHKlU6uAbkYTAKk2QZzLQq0DPfYNDUyLaZKRjZ
2JvhC4TIk/7o3aUWHrg0HPbRD2L9jsjEOjiSdROfcHshhTYvHglv1nxKYGfFOlirFxwN8XDO9NQ/
l3l/DamlKH3Vk0pC9kgGx6o8xeDxZ/lhjnzWN/nOs4VrFpsWxNF+Cj10MgEd8EMkp9VMtqjHBJXY
Bjiw1j1G+mB2YCJZ3Tl2zSWoraqLUt8c/UIMZO3AoSkCb9z5+fQv+7uK895yTmXPcas0uiVQbEi2
QYdIWeCnB0LYA/alY5E8AHAlmEgmZhOQls65SZJNL8v+xlwB4z5UGeaLQWtyftmwHgY1FFYtRsGd
lsrZSQUuDXa6+xoKtIkWwmlNJi1D39/S4TLRKP8W6vmZrEFc5DxQ0fVVciY3151Oigq2sOYJOPhk
6sAxcyYiTFwKUzeZeuuRk6CoIFpT1g8IipZRfRYkIIO4SMjyxsdhdMurjjcFm7IkTAvyRXuadQLF
8OL3szGAS6Y5e/KSDmWIk4pKp73DsOrTp0jhG/Oy9UpDipSnnTboWdjeM7/yi0kVsyyrhxIA5oeq
FI6M2/iYUSEv8IEctJ84rj2BDesrlxLK8H81wKx0SyEXBGEGARioRJ6dWdrJI/09rhVnd1KO78B2
wTaeIwIeuI/gw0dxNca32MnhFyA45q+zBdLdrZdQYHM4E9QSKWpOMwQI5QKNH5xm7Lgb6Q1NooOh
w7aWo0/278NPByeyvH6dWthmwcRnY2vtWkt9SdJxAPbh9Gav5IRYOj50yUbcOZSlpQ+PoVKTl0dd
A0rZeQ/nyDvZ9MhvqbmVPIXMSfRHBZGQdKJ0cjxHFfct/xK9W+kq77TeEhkdGhU82uc3yZGs0w3V
zo7cNo9H6A7W2udHD7qOY3PdjDPDyKl7bbUb55v/oryaOPRGEJJu/sTn3IXW/psfWMdswTxLRvTL
Jz/R0APTLcEMZKGtVuls+V1cjv7BD7e1G6mfxb9hDVtQZOc1j8KW2GnCF5/M987B4jT0UywlND3u
Rma+Xwo4aP7EPPaCl+P52SQCHPJWMWyyueM0t1ZxeZANVzxMomsInouVn3amJXh+QlllAA2uupwc
E2Y+6VlMr4VkeNN2DmadUt414kohDc+e1uTiadBt9XmQRuQypU+ipqugqCozCbcYORqwZAMUHHFe
tQ+V3Mpa/Utr/guB1kgjio0VTRH/pjW/mNbyl8tdnFN7msrtTaJt9UJYSmoqYpYINilGurpR7UPA
pUrh6Mw51MJRNkdujIrlWjUt36ELuUygTl54oowaOEg1Eo2BDJBnCFk57fG6Sp1zeB5CeEWM7CoN
xJZqFgiJUa9jCCbg8ThTikjXN+8BA4Nq70QgjYquDlSsfgOOWpam1kJEHvbvZPp24TTUWPkYgLLu
+8fLatfa8WVgfLGLCOEpGiCR4edDx+eiBt7X7HqdCynewNaiyXKH1Zm/MEB6+LZbYrCLUfXtvy9y
2YG/Ntl54TMOPViWdzyxuLjMp/0p/MgKQF55V9OhqnkWx9o7AuRfuUgWrfwKAjbG84Y69+kGdNzc
Pi8KeNr3WT/Yt0FD+NCswxXS0WgH+6pP9PbtdEzqYq36kXFZhbm19QYcGTLC0ODv5Kp1REURZINZ
RCVlmNhiwdZRATqHDxpXrHTH3y88IRQv1sZd1QHcpISJ4XvJq3uu22a3wGPrmgs6skY0msa/qrU8
e1G1JWi/94cDkcX/QgQN2P9QNOoK8OMncwkFtDl3t0VCdNOUqg0xXK06Lq6UkTUEohNBfTzFbDyG
ri8huDbGFYoHi6yOV0XmCBCwcR7j07mWl9UC33rQoxgxygK9YeS/Fxkk7O5e4/bumHU5nzAZNAX0
s9rrrgw1agFTMDfyKHhtFVW+ddThLVhliGgc8llwSBEc6vSvCxoVbQT3gFtsiXKUITIyS0UAb7tU
kdea5e6/KQJhQ+MrYnk0Se86+jg3C0RfMJ6F7LAxuBpLV67EqUnl+fz6/X76G8kbVkP4txBWrevt
NrmwB9KtTGlie8J2X9HcSeK4ZoGBH5iuCfmn2r0vNS5p6WJn3SqHDt44W02MtHReHakZbsjMKZz5
OzItxbWp1NmThMn2ep4cON6uoTV81pAUJkJcovh07IgsZWMpJRC8l+5uut9GZtgLibAAPWoG0s2e
oTSpzQ9732t9DVvJdeSR1CsUX+JTPXSz11X8TsEHc4OCCBY7i9jewBuLbexFYHPJ5uvzMDDNxUls
aoitJFkZPbx5R41DN5i+qeEj41K20DA39w5/XG5PHtr/Eenb5m33LAXMIWqnZvebyttJ7yPGNrpW
Ug0bdG2MUbQAgBd9mwCzDpP4jp3yMHRUdZ2u2yOmADxNGqn/lGWTiWoCcyVjDTbXv4ghYHYD6y/U
QA+3n1wGleunyCK+OYM4b9T4FfYUqtV9rmzKKe8IYhb4GFlh/y0jVxOjXAH+cgI0wxYxTqmJuPkP
TT4htv8ZGHCXjm4GvcgYd061EP2G8NTX11hcFzwxMFNbu5ANwTkMgRlLlBJ77HGI46qnbWUpc6OZ
OvZW5mXvGuqkbgPrm1LZhIcpzJbwx2TVQNgCxE91hktUknTBhKGxUkp5cjwUj4V1tv9plFdcx0hi
njxd094mYPvTCsVBBF5ANlReTZMVn/y3CaYr00B0gs8Mqj86kYYGdjEVr30Q0axdrIeq9sklFa+4
SKD3a3s7FkFklMQylctHx9RQe+N4VMfNeaq/R+37vKyUgot8vAexqYXAyfFFDyCD72QH4xRz4UIi
Di6n0CqXaBV4qJv21rNL+5YHxEW34+a2y9KocbbAerZAXhgsXRAUPdEjaoTLkCd3YCg9BC5I/vQq
zBJ1HKXzFlY8tNSDJBkerPWK5GO2iBRbjRWaKFaG4fmemMxygo/OvGpWsgL+ykKMRmuXDffCqIsH
A1xv7RI1ZUy9Cwj3dVWlYp3YEnJgAETe4M9izqcpAiWnuT526xNUjGR8cNF+3XqtoWJpgUDCB3Mo
CRqtfa4hP1FdrMJ+KUzpTaySKzA0CowbJSjQkraXrsuCoB7Cjchk9m2G1p50qecs+eM1qFhzlPFu
zPtvyqmQzCGwbfmcTzOQWcvgxyKJrweIp80ewxczBMtmJwega9BdqZf3fuzY+vw3CShW3Jh1T4cB
WFXHmVNCxCHfrTmyU0A8MQQg/CzTl+McG0No0fiqRmUH5YpAKrDFxpg1J+gpCDUYrSu4ezIaGRk2
w5tQPoKHQ75nWfhs9tjZgG3UrmrPhduuCHgNeux/AzYP5gaHgluZ9rsK3B2zS738RyR1Fl/NK0Ll
AmChXn9IzaEs9ZENwWw1jSWwe9HcPhEtpFwRpez9W4bv+s+ho9KhINECCm2Gy63EGktbaPGHvFen
oCbEhKbQNPdttwjpfxeKWeVHqWNGNmoxGkUzihicCevXLuyP7mA7czuppR7AlwE0LN8g+jBJ+uhT
Z+1IqrkWMMDKXobPGGaHLLzeT0RxzNlW3jGx8NmBSvEXNxCM4s1gHJF0QG1nS+uM3Wl0nYmjJM8Y
z8sH691hUbMYry0Z48KmHruPEu/RR/i4HeO4ptw1elqVrZJysEPXJ0AjlyvUiYW4y5+F6mGiGaCT
vaw+7+V5v//R0ENzv45J7dtYz/ebjWjyfjuK9qsb5Z8LeFo2s3eaWl/tg6LqfjG3MCksT5/a3F37
Rm5lRxL0UmnU+hjsuHgYtkEq8IxunOjs+xwaSZOnoVFD2XJdeYdtmW3RUroO/hKr9zFb25yjkTkG
r35qfUAW2+Q8rHqdizfdrsG4B/GVSnyVZYkGLFLL1Klkg7pwQGtnJuMvoDhSx2gFmNbnAT06OPhn
6IK814XSlk2VkKgZYvu1FC5HeSIBMkIIVz7y1fRj80mlNK+tazG3O212yzLE4WGZwhe3I2FU317G
iAJGMwag6aQysLqfGxtMVYpccTNgylO0RnF4QgWurSm539VE1gh8ebazPTfhtkb4+BkYhW5dLTcf
tuVUz3upVtQ6fL+XPWWqr2AgSMKk6Hto9fu9Eo/sAEFNpnTQNUPyGMCsjFhWcYVkH8V9ighu48ko
BqYsMVg5cDirM1ZAB7UQ9NruvR2KZwZiHrqmI0OAuUXybHfKBATV7IoytnSB83+mJwSCaG6K00FP
ZecI5C20gTM2qg1kPEyGYrxLlR6xWPAmN2GNFgl3yKLzH7gRUpT7VSshkpVpx2anUUIuSMhcBLzI
1OpnprICjaxSHGX7Ba/rVaRMTdLK3KtEmKqFDAxoK13QZt7QJ5n/qh0aQtVUKhNizpJFEdHzRoyB
7ORWOeGp9t3LM77b0YLCaM3MDeD9uUiHVkPKO2RPSV5a7ECbpeUxWu1Ut7tvtei20gUx1hJE/3dD
Lv/uD1RnzVxxlVtKbDnQD+SGb4vUBRfok8ceKm03VxvbuPwPqeARqyjZ7BnfIHJd7a1OnEJy082Z
rcysMBAADFutBxPAWUYmeK2fy4RFan3Ef91FBrJ4V81tuMQqZE7ecP0lzKlOLZexJ37rpiJrfC+z
zlNLcSbEoIeTry8qCA93emNu6T4FcuxphB9EKeT2alm6s8EpjEgDzOmh18T8xJiL97rtrUE51YIs
ICZ9vPcLLbB6dp73O4BUy2k1V3o6t8HjWb16M9xnm1pZ+xgLdYpI+L78DdgjFz+hbxh3piUyYd0z
xiZCsvyLo1NFYcBr0l+IgGYxXrBjklcVSHYM00XvmK2pMRJCYoDZjpppvFIBjxMABjrGZkdQTpTu
73pvKyQsckBACt3p92QxEppYlsCy7H6TxI2r0vnebDafQOtLbqX8kOlK6OMde+HUq4Y0fWilAh4h
WNM8qnGwk0D1CyJVjr01SESVmmd+MA9HuYOaL5u1XjJvNIdPhMZb0LjBUyoyLaJGmkpLiTL3jPH2
5pSZc0ar0sM4MecOTzfM1m4hMMQcCNRmZSRXTyeBp4Z7WR7pMnF3v5BdYtn68u737RJl0sLrBkXH
99ENRo7O1VauCllrxwvKMzON4SihvGEs8+hcGLOysiYMEXUi+bzM1j7yAYylHwnJQGFFoAf/kD/g
tjsaVpBwkZcrDo9g/EgtYDuITwgceBVYpyyFIdJyu79aCEr/ijXqU+OJspnGA16YNoU9eDayiw15
ZnGPsoGPE5ncdkcsCS17Cm/tmcBIf0u8wPpec9MvAy7txONcraY+z18arEnMZegMH/Et9S43lseH
I+R6jMrUMLmEmLFa0r0PkQlhH9mwnTSw5NAkuh4xB1qPRy41v3EYqeivPAHyL9l9UF3Z++qxrWd/
0ipQMPIos3aQis7rXcssN9qjXF7e0+X3sUHwQmLOAc32e+mECtaDwrd16D4aL1rvwIopVOFS0+43
P6t5vhbZ6vQvxINf06VH69jxgr6EolNMTQzsBcNjexvJgAMB5qHUyKCeWpc4u053bbfDVPnxjpGf
nY6NAIAgLbpclZJTFhYb3Rj0fiDOu4mwy9BNpTmlfWucTCP395QA0sQuEGCc0F1yGUB8IPud0kEG
2bZaA4mWr3EGRY0o+lftGAaAv7RqW0yhVt41uxamhnpzTtGVKu3WykOkBEJln8kbfdDLGW+GbAOh
alLQQJi7ZyNcEZiRwpXNQMJ8s1k4eyrEusQUdlDd+kPAnDLO/rD6eWetzOfOyVMMaRtR2Aypm88o
ky7sZ6r0MONds4TXhWQo3DG56CqxnHClgAgFBEvReF1DxAiy9kYV55tOnRcFyg/PTFWDd9n0ympM
PyRwKpj01kIFKsDgRt0fNd9KvGemffo00aazeHLVs7OAr2rqIjiU2kniwCHdFASeROW1dXiT5RpV
jkd3F7VgXKJ+GypOPln2rV2b8tN+RngcbDfvGqFxj7EEF1OjSFS3bCkUyTP0LCITSFF4lFPRoXKU
mzoaFTnYBWT2nwRpkn8Uu9AA6RWT4txpDlRfkS2ASgBe/7+GmBmBlIMHkg3s/rPoxrEFBlhH9QcI
nyTo2zi2+QrT7lyzxSHpLZVMwZ5MAE/pUyFJEwDNOXE9x8Oi+X94xsfjCJa8glFQw4hx3lelztAY
sXzLBYOKqFJX29/HCV6YQTcuizWBbO6ueCtNVmM5doQrzO5+aIcrJiAZp5mWFnmcK8RQ5xtGi885
Hjj1zEe4RznGlEnxYUrhI+BNNYp1aZnyZjgzeLDK3wgA8YGCp5Gto+GgD343kIVY6xfSI0DpuQ1c
tfamo8r9xCL02OHwiwWD4kIgVSTa1fqopC2O7gSFHAppIyJE4R5CttkexXjGOgIKPPoMNfidHrln
2r2QxP7977irFnblV8sF6ELc7TshnW8UMXo3lHYa4Nz2IRcMs6x5lPyX5IlVm3nFTGFyUtTNb280
HfKOt3FIeG8i22ITv9AkGxv2HYXyAHMhpebcutNcq4yL6+RStOhCqX/gk4GoSFWbW76SxskG/7Qe
svDKMTvvzodc/RnmDRvinhrmlgVs945qn3eaf5sgzLXMntjQyCTthYCK8GU4T1MZa+V3U0DBVtfg
hY23DeQsdKvfYKfzHTa1BZgo3sVYtgEtz8UyfXCjFBFKmDdriwNZleUX7uT8nQe8VHVndA2wjMn8
ONnbW1ga2NW7M2QRnc9w8JwiSaiMiroMnFwGLs0mDijYJu2ejW/P9uvZIqByOzEOyujKBE1ORLKA
5RyteJn2svjogl6YawU98zA6kP5BFX3lpPI+msJyrAgrHd5X6G0PjKrZPj8d6E6Y8UBjUYcTJeQJ
Z2nA+oS79InqKoN6fZOTgvLnVTV+QjhSIkbCz0o5GFFQ9VXjp6e6XhqGvFeki3GF/HVIi6cX54bq
1CAVALHsZHvH30xVK96OYpWOHxD8OaI56XNcrmfwkMoqABc2r0wqkuhkKDrmB4yUBbaBJnP1YMUn
O04kXWSFz3sh7cXLzMK/2Ad7RwA5dow81/UdgDbTGhKgIvZE7Uo4WTYqYmdkUN9QYrqYdzF3HMAU
CrPbi+OI+UAAi8aQtpCGgiMngvkljLvObs+OnCOOAssOWa26BHHdPDYiP8/NAjSN2WGIxQfiSH6N
C21/o/zOMdrM/Wh3OxOhsQe35U/mqG0uuz2OWQP6sjDCRQu1nX12Iv2bPcL2inl4Jp5A4wOEL80T
DYeBQeUxZoTqq8LiNswCBHj5K5tGFoccwU0JknbRettz3a16VmQHGr/iDbk5bnq+scppjPGxDuUw
6hgbwGmBO4oU9MRqMz9DpADcJF45e0hlwYWuv7gvBQD1cZOlBCiCPrHSnGFv4Gv3r+bp0p5/ROMD
0RtcxbPXg2/ARovwqUZqbixP1ZLLho0NcrfJcf0900TEiYJc6HWSOg3ZjNCZOfs7ALnyneUShryF
ELY3frMnS6kkoNlgU8E6UoVOy03Yc6Y2bxG2A26quBrKF5AQiBpU+zhOLNfyso3FNGBM7Hf+S1oj
+u0N6t9QwchepQ760e4Q+LI1RXwTWa7UyaU9F0aFhmMMd52Pjk9d6vfpi/2l+GeaM1pC231WiDeK
8r55gd9Oh0U5iY4n/k343mxLYSTCtKpj4mYhPZpLLpDoQZv3Mno1PsWH2RHSOhcm0KqZr86USY50
hLwyklLmJhVQL/ImoWPjtdjmE9BEPrCG4wRrM2pRDrpRGgPo76ozbYJujZQ7U+FcROrY/hbhWy7Z
pbdNhbXRXOSYW7TXzb9LVDEDhBC/hig+quMbl4Z4xt2Ik8kEg1Ev8epW+zS1EMlMP0kon2QsYgNg
kL1sdQLF2J3XP2ELWJKefCwXW7aVDh8Zr+W2XiagoCkdBIURDmny1EZYiCOWotIiB8d6b8rVce2x
rXO37dFKtdyfLAYMY3ufjkSgzrav/ExbAUOEYlG6U01QY0s7PPhJTqpbfL6uhJf2L6hik5X62p+G
Xy8LhsMIF9e5Szhgarq/0qtMEFjd4WnwIFhon8HPArRhVRhI1VpivbrdjN5ZnHh9YrattQoZOA3O
K/JmTWJe2QaAgf54DKcbVy1PADAhtmW4arrHOoea8hQ4DM1/2oncl9vnyNWx0cQYPUTAR28+RJ/K
atA1aojutbhSMD4WUCbFICAlEpYM9Awd0YNEi5FiMoKai1xqZg+VSjg3b/ButJj9ABA5Si/AzZQ4
DHev362lA56sQ+1gH/ZWzekmYOWCtAuNLYtex+LXvIURcm2pNqDej+Zzo2wUaWFY5O3lngPD0dqs
Cd79dw4EFFScjS7FobcBfl5IHumfQwn+w7Drnl9RyBc2ff2U3WaiATMfv6xIxd7beXdmltrLBfFj
D6m6akAgCfXOogppfuUb5Gcnglw6DALqae/4VBsf7oRnXQUpcpS1vWsACqZj7miTz0vEIF+1BOAQ
Bh8zl3qONXBJ8U37vvZ9Wm21VPcJ2HEJw5TOGfzG7VUD/qTvvLn5aQRfROh+gOkL4zPODPBKKYWN
hREHV11nkcxiPMchiy0KXHUXiCqIG8gTRj89EPJ6MAcodK46cIu0maMayOjhKtXMO6qnTJnKvTfU
SRNMzUnPSlpC2iLI6YSjjg9Trjkyh4FJ+64UKCgW+xudtcOWcJ4nRjUphp5YmpUNbwigBNSGfHQo
1fYkjxY34kTFo680iMeeOabXCxU1hgwcKkc1mNlLXn4YlF2PFTrEK6kxrWRmpgQ9NGhScSdzbyks
8KVuFFLRQMUMbsWi0Jvd0+lFNJcqYc7kPMghcKLnw+4hIJj1J0EOQjPHeN2xBZTgMv7pC/Xs6gUN
onEoRMbe1SPCn/x6dAiTW4mbS8pAjBHLrWFD93ACdpCRLHcyYY7KE4pLa1C4gdK6Zmw4HsbQOdkS
iRVWPYmJCbc221rpJM/AkXr4ocHbxwxFstD8gJ8yiTNg5nCt70sPuKtDPgNyFuF5u0XmyuWQ384g
al7SRJHEdF+b4/JGY2e/zm2BlgvYvutju6Hv57nCPGdeXJrVy3Q/hFVU7K5pJ7FymORzndfBMnb3
DmLlfr4vo5n8kr36GHrBmW8LuEf3mOo+Hv5f46PTLMOPFcU2gpVxd9qok6Ew/vLfKE8/SBWKdMB+
e0CoP9G4XHWRHxqLVtUBA+dHTWRv3PHuD3VgWjngb4ZZVivYdX6n9o6AkBZqQOV1gxZZ9qWJiocE
trcZ9uxTYxSsO2mdysX84esh/a1JYXiI2FjVOhufz93LmlnS3TE2/CRoRlkUr1aujjxMpPOoK/hA
Z66JJm8HOoDlQ3YRPt2Sph6ew3RjEkH8LZjnqCH7rUFOLrfc6SSMRxpFECVc2A5jPnNHSv8C3Av4
SuDA4MiFtAsZvOwOMlgWUiFbQYMmFEI4CMXDXczErH3VczmVshtnSu/HAN2jYKMi5cXVAeHYISvI
Xdbaes34QJDeyTvANroA3HENQwPBWBMg0Mgv4JJ4WFYJI5MQCpgMadagYtIMihXNYXPekWeUB3aT
fwEVg+LnxfH/glJWbWsBdpxMRLhyRceE8+Ai1DrZsCLjzxxdR1HhcOxjvaa2m2pGDSgYT+jDKlKS
wM+qvtwOprw46Y+rxjpgVSBf0JEu+14H/ufI+IoNZuaEpUfz9pB6f5KQCJ1yg3WVbHPi9Pl+wTL4
iTgAyXVU/17IxJIODKCmfi7IKYhhhJY9PqkI79PXhDLDbKgNK3WT2kq/HDtG2UWMfNSX5cL3DsN8
MCZSMd3PLIQiEXv4elEYEMfypBAkzryIzlbaXjCQKnLIGUrFPGbrX8xLReZMieVI08X3S3pZlhDX
RfA+S7etza5iNZrS4MVcToKuO1Vibhga7GiH2ea02ncOS/Ewm0m5SN39Vh7QOSii5BOGJKN+SYKG
+1Fi4M4FZ4DANrFuzQ1nUa6ZAEXj3h7GPH7mDA1GQ9nCW4q+XT00pfKa8VyTbE2AxlwmH3e5BkCV
rNmND1INiWPyB75axwZ9MS4nWry8GbPD+F8bJ8tq0OOOyR2F7uKc7x7xPGZW5OgeLRYTKy3e3Nv2
NslfJHEXE+dEG2FunvYdogTcvgpll5Y4F/8XzBqCe7rW8jx/cOmFWqopl865s7SNm/XPZ6wHrKWL
LACS7kMkuHpx9KjvQ4wlQVbLv+qJNk7lnaQpMX02dw8+PYXnFHNU+TucYMZZHZonEM36BZctiZe0
fAZO/c6hdEcHvZwIg2uvW4A/4CdYYDU8JtX5IZ4IMn/eZZoD09DeRDJy4CwF5YzdaYB2ucThttDX
A3LLZNT+bDkJmSH4ZgMKDhE9RGFNSnpbkvg8LD83Nqiz/HMkabm+0oE0A2REOP3/jio92Uxt/jvY
n2WfZ0/bQSKZ6y+pZkx3E3txFwbvt0i5Y1k9mmIuzdh7SNCKulf99lCNGBC78LdxMOx9keB6KqHu
SA9ur2vu8yMYBt1COsNvVq96AEuLV8gZXp5CJ1J18E7IKopsXwB6Sddv5Vj+eXQNaIOWBlsZtxNf
au2uyTs5kPM5LZ6XgaIPZd5LmXv2CGVG7KZCOQtLRS4buiWVlPJTUTqZSmspea6rgVSvctn4A0l7
zYnzoRrj2CuyEHK19bxPs6390Ps1+Adf+pNLKeSXA9OK82nislYFvZYTFvSNpzIlVj4/rV7KKuCF
m2NzLcY42gLtcPHq7zExkEnAFyECtFI4w2RiPIvExtAYM6Wao4fvZ2W4SDjdvcXylF2tZfre7vtP
8ULDRuz7CJZbFLFGy5GueXeIG4kXojeTHYY1BZx0cUeLrKz2kZUzaWh9s+k139DxznYZSqI/0NPz
b3jnHoaF+SzDaIaptCwVziDUKt0bzMKHFvv2sSZYsJJeAl/pEXKIznJfle0hkFwyip/LIv/3UnYI
eWaKJswaJo6JOCioOkycalJI5RDlrFL4n1SUg922ajf21XA5d2bRcGJsy8ZgO2yPgeSUqQcNS2a7
WiEBMEyoqe9tFgApU0thOWgxpRY7mBw8voT3uroE4IEYCdj/VJxN4CJ7i7knAsQTYqCLD+5+XtZX
IFhV2Ko8e2PBZtpLlP3n54mYQf1FBsnNIa/6uPNIPwaU9c/wUICgNF8cUPf2WY9wYBtZdg+SQp76
BXEId7cJ89FXVN8LWTbbBNGLyADZGlveeepwmFx+2CalXKWHniJR0PlqyGg2n02EUWxI7gDpmR7X
MZiVmtxUqVW0FsyHUJneQpnFr8u+hq2eyT+VWOV1TagKIaxqDI9D0cKemI6XhYvy2lfvVu8aHCn5
Zy2iGjHRQJu/4/Lcs/qS/lN2eJhWbLIznpHe9Fc3SprYdmEUGVYgQGAn4XaLLevyzNqOcUoOc8q/
aPtE1/zEnEezJ2C0ZCy0/4cnjZP9q5SbKBisFIbYyGoXUCWKeTu67X0J97IlGxHO+kbl5Z8DBuWt
w6f0uJ11XAfcjnzXs0ELZGoUz0oUm27WhGHlhQvLQNsVLoGbfaXlO+/6OBJ3VOu6u0aOLp1YgBJI
R1/hVBMhRsfPLhVRW5BevZ5SEtE1nrSIZtZX3ziJMBXOzaBu5JMVJS8y9Fw+ptOYzx2PIWKpzW46
1brpT+UGHxEyhclB0DTIdqPCDkMZEeIioPfDTxViHlx/ibp11PwvgVPpEobudChi61i8unRFVVG4
0btIumpwyFwGvWSUmoAt6KQKRkQZ1wrLXujvK0EthhNbNbB89sOJxGCdGGe+6K70uR7WHPRjPqS9
jwX9cy+NK/feN10WmGkkE+11+V26/oF85RAqAJJ7ecLxy8IITX7z1STXCZ738qv+IsG6YunjQ6ft
x6s9u9rr+3HfauPPF3eDMLnne8pZ4XSlCpr4z1hC6PGVftgbYmYmvqUDcHI2wyvLGn3m2It1sN6H
YqG6GrbsUxEBHc2UNAp0rFGcA0t1Z6ALEOqiQeBxduExTpw+eZ/Luu5DoXpP2s1Rch8b9WlsI/Co
HhDX5ITTsHIjGUr7XXFWaqJBEoHSfkHDqSNHJ/+uoUz4FmKWGA/NIj+3+ZtbpRj0lOMIzKmLQEmC
kIppD4WgIkdQxuub+WEpoDxETybhraWVceC+5Pnk+IxUpEExV2a40+xVzgwgNav5usP8FDAUd0XZ
IhzUdlm22R8UnBzj8yQCimhaFAo8nQ5YNEffFAJOGyeaRUGvdwRUoNoJ6azDBl2brJsCJa/YF4nD
0EwXfkFSEXW5unu4Jt4it6M3Nlsj3u8u0L/zZ1Lhml/RhGrwPgt+xUmhBgBinsAmSd6xzq5PxKS/
ZxN4nTNtIXIkTJAAun3TTlGxHzER4QfxKQKRqnqurKp9bTzVTnjkQtgn6a21vnAxuUuwSNXde8+w
wL7uLI2Rf06F3di3Ah1yVaYdMSFVpEMYo014VdnjLIPgYMW0QQVsg1c5mVUBI4vxl+1JcRcINUid
kiWOa70AeFM7qZj7gOTvaMgMB73cDkjrPIc8djKT4He2UY8UvXxqlxGIn6n4VlsFalsT0O9HMyzs
fL3OKQ1q61nP0moE/9JpwCYH7ga6Jgrwf4/0a0SmpXKz0KjMzgC15ZjEaWZjdBsHnxnKsaSa12W1
NGUWA/lXyQ+tQvrE4Z6E9pFCPl0iF6F3gm3YXLKNj0t9Gi5RZH/7eOwx+CVOLyAaDCXaOG7TYtV7
Q0x0smXi3g5wtxR6PtALVMCmv5iXG7jcb0ER7p79O7tXTaVV/YxoRDbOYCNxu6mYiHKAqJr7nWa0
3sAcX75VLBYWmpzUbvHveEjbzI/mU8A6WEXilLhK3AGfOGCx4+7ugnIN1o89QVk6ItAOyXt77h1Q
9EvidxKTy5BlZu5J4MxPi8B7r3WCx0lmypR3RsEbjIRxFQ6Tvx8FddQhcO+hx9pkuu+wbNYjHEFm
UzoyL21/pItWIg3uDworIYPJZ2uH6RsnvzJjI2/FcEzYOW3G9wXsJuVMFeX0dpIrGD6sXUtuVq1S
PecTb3PEHudbakGdEUnQ/KvjTxSpSQNUxyz2F+mmcBI5E+Pri4vc9z2HXyid2RRb3jqquywMZWoc
4x/ZJ/dVko1FPQmukOKyEwnYIer8A0sLy3ZYb13pKeLLeuz8eEW2fAlsM8/c9kKil84FhYdcQmDb
qxHVU01AJOKfqBElB+8AnucX3TbxXhRLc2i8KiXDK27VGZgu6grDpQu6oX8hXCTP1ZpGIvFgVlbW
tkXGbZFEdhdmLzU64Vn3JB7fy3D4Z2dyf5EBJQjNV49XYeiRD9PO9yBI4X4KeRnPEBFyHD2ZvdXP
yEt1bn32AZpE+pi92d8MirxCe8orEBECipUnBHcBJnjm2XzZt6IeW4ob3hfMAduJCi2zZRImh874
eDzrhjACt0DnwO5QcuORShHQAXwct4fCY+Z3wFqWcayFWtGbYrLCRly2v0J5dTofUXBEpoM/nDMw
ztEQUm1IqNFMOFozf5kH83S6zYUB4P4tJTfABxJInMfFzm61VYoYeUiyKWatuv+mszzqc5YxiBVL
vJy0XMGGSqQ67urUF00Pq1sBEUTUb930150Bl22bJOwPKpfMci8VsuKjgHIycnEwBvUU+NlGBlya
frnGSyTbaSA3TRmsVoLai/0UT8pWr4e+7byDkTyVg3C62a62kOzPixBwWbjxxmvzzXLAL4TI2nU1
l7SDK4JGICDF9C0VCcOK9ZYw/av8cjeyYt2J96tELfoVcGmqpKVouh827furAUEipVprxTm4J8/W
+Tl+Hd1L9KK6pfi/FysieHSlp9hMDTcr+uPfKAuwumt48NF1R7kqrTl8xQTfzBlMkjpkITJ3S46Q
1QY4NhcZRKw/Kq2+ADKcWYnI4hkvi8HFJM+++3VQwGzvuMuDzw1LM9B93j0gpURQfbGh+6vpfMV4
9QC4caBol8c9cUIWOklmn3fG6e6VXAIq0ADYbkeZFWpuXEQ1M4lMiXMkriG0msmZXXn3p1qPFvou
nROVXDIitJO739yCzCAToRDCcpti3Oaq2rMKnz8Ejlm8YWE5aHrx+iuVcUzy7LQa+0koYbdq9IWf
Yvh2M3FBocjNepCjHraI0nMioz38Y9XbePQFWsFiCR8k2lYuGn9r+07oyD7kJHW1YHOq+qSWk0n5
yPBAKTAC4c1P9Ngdag5tWpr0VxUgUaeEivFizm2r8YhHGHOGWL8IWKgj8KChSiN6RRkLUxM/fPse
D6KX8EwXmwkF7xMWrAhhvgSpBe2IoUZxsrqq8+Ex0oJRILWE+en2c0oefVlNVAMhtNLZmlETdEV4
GmzrM+e//fyqc8LFWQWHgJ8MWD2PdyyHKwHWbWswfAErRWIabyiN5ExaTQPY+pxEyZQQFhJ06J2C
d8I1xooJqb/1YLKTpITdXywcbwYDBTG2ip7FRVdwVvm617GriFVScCjG2npbmW3EzESr/IW3IEEf
MvjiGJNFuo18GwdWriiuBbTDVRLmqB+0LRZFeUkfRXUpVqDEPGNF7JNJ6EruTG5EAR9wtRZbvLHu
/3BeND5cJrNREDcBV2gPxPD6r/mvvYrJ4un99arWdBZ8XilrbfY+soJjtZOaW7KJB07uEREVK1fy
Ymo5rGSzRRTAp7lLawZWJpIWTpSVSD1cp12VOA77CK4zjN9s6Jh8Lt+3hYvT6jAnhsFwUe4bvEsf
er4NgB1duQytSdIi//n4cqZbl37jY81RI1r6FrD+vODFGw5AVxGlvOcPs0fjRwgSh9fJKHvoeuzW
kh9iGYpWj+zWi9TIcVNkdD6GjJYthkKeWL9kCrKZTHrMa8K4misFRJ3kIOy9Lm3MmC4jRM7ZvxpH
aijUwQ/kenJGQdlDnQeI91s/eJutQfa+6pHIq4gSLlbXlMAAgxO9QCkcLJ6bj4lau1eZ7UoqgYKI
HWiVALyJoMWzWg+wpIcMsqoFcO2XU/NXStv5vbLh4FnwRTiRL/Bdm06g3JXx/C9w5aIasGMQ+1bi
cSpTOgIa07lrdkuGcQGINPcyLKJk5zoqTwpFD26jHZAKWFg1vqyYYWtluq8dmo6qn8KlEHsRU7RP
2L8sWN/ogxMfxuTu768ojcDovGUjZE7mNs2oLYefSuDyjx9Ri9vVS1uFgojD5pNenhcmo8CIqLS/
6nuodu2mvGWmVv01vcRtaUmi4ZcKX/2uYLkVNPY5ojjyiZVJzDNEa4Aw+NStgoeJ+frYtbWFXhmI
rgUhf1NLqkFPdQoyaqMr4q4jYkh2RHqRtQ8V8hbLR/83Tk3ME42nalSZmjbi13ocLwyQiBkkzv0W
D91s8xkcaA6ChQMU6i92DzcNxTrXIcucNsi7URg8hBLsLjqPZ5TBQSjiKA3F60o8auCBD0N56TXC
efPj7oPdB/cxRaxD/7YcMVzqd2EkRFRwQem0grj1TsmdSBSfQoOTdywjj8koEB5k+MCcU/jMliZz
1o5nq9p9O4ruWxKACUennGYMBLD4JJYdM+3ZqvyTWjIsGXmRzF5vBA5xfjqNKf0eaKPgtTrlkBwP
OjroeSjkN+1bKjbOyyVXAR3lpwi5sZyISDuQk5WvV/UtZnW8SJdu+HSHdnt5RJFhcBXE/WKUDsNh
viz2wg6aOGSdBahokzWmfI0cpGvGDIRfhiJMVuOPMqKZzez0THVEGaqT28k0PebgGkPWqLTiwcE2
QBYSVPSPi+ixQ89IcwdkhI89NUvFuk22kXZD8P+7ifVPACpCNGlAiPJnG7SFPF6582yggcK26Tsf
wo3j/Nt6IkgiHFLQ0geJgKpEZjeeGfsfW/Y150u5NS35BZhqRj2a7wltqJQFa5ulY69KwPZeXE8q
mvLgGyhlXDKFRP4ObaiYyuBe5AMajQVzxiuSJRAp60f4gPBi7ZOIMK3IZ9Sryt8LUsZAG1wZUp8r
ZKLy4iNM7WO1MT7lWIriwq0wVoRt7gdOpDdVONoSKzMUd/V1ROBZ7k7E7N6s1MAwIad1kJSWVuAS
5h4HX8GPQOmXeLERt8UPcPJjuznlRwHxoQdFP5fzXpnD9biRFvl60kK2C/U434IlugnOh1Dp7jQh
/PiFSanxcRmcs0G0zVKWHu+A+wv8mBR50uEl07McfhOVMSgKbr9L4RDATfkKZ4Zm7Sf7BcndAAXJ
1+Ri5ihDR/pECwJEw8QhSbR+C48UwZ0pygbDpjZnMpQjchV5ngZm1oxCRfNqHeoqDFke7fOfMi4A
ZfcjZzABseuGr4lw7lnqxZmkeBJz6i/AU8wGByqHhFr1xr+MaCbKZHNg3kLJrvAWmWJIYd6e/4GR
S3Dq8lglUNtyjFEEOlQYEmitRQd3yMQ5Nm9VoELZkf6TT3phX7Jd9+5lpwj8LFYYX5R08vVvVc49
560h0KN3fPPJbyq05AYQ7ZIVHUzFTBCmYGyPY380xj2ZKI9pa5uasZIH8OL3sG3IdXnPIvsvCowQ
2yUH5GjowHfjsBoL/2aSlxtL/sMpBn/YDSfusISKJ1/hrdjnf8AFhYh6mgDMyXPqEDNbjUelSiaZ
mXUo/wyuJVE77LqT/dKU9VkjrrTjcxIvcuZpLw8SyJ8QlMebzMnvhQff0JKc5E0C4Ij8CY7KXhuS
638YpQ9IYYk9dN3RezxxsWGT1uTyaH20b/gjt08te51638zb6CE8H+BL9eI4YmJY30iAZFKMAGno
iI7bNPb9ug34N8focdpLKeHmF4uI0qks/SNISto7uUKlgh3npL6FO/yT5XKx4p1YQWD/BDsq4ZMx
P+mwqMf+wHXdN/iKsXK5UH6MKyV/4V4K85zwY7XuZd/oou3OjQmGB4gNK99xfwyUihUTJIR8KyGU
CuP0eiGJdMzGL9ho1d0G72BTsvZlNUXS9oiw8YQK0+AmNiXwTNLtcBR06v5FIoyrWM19eSWVrrN3
dXoNLD/OhKfmhaIqq32jiPb3di1hqeKKoBV3sJtRmzKz53rVrH6XmO5ex988MDHfT4gjP+y5VoDX
ABIt4L5dFde68BZMRoS/cxl9jwCWTG0RVvOOR3G4GvKKIPU7X5V7u8DciVeTPY6JlWSkt/nvIv8R
zW1hvi0RfJ57F9kmEH/0eI+uyDZhmj/zQ8ocPi3atDlZ+RwmpIA930Ect/2tsYWDb9pTg2r3wnLS
qc/3D2uZhxkwnYYKz0C09rfYIqf4d/XT6snStjgDSsJK4tyw1WgIM5H4m2jr68m6L4grb7WhHb1n
f6UIxyEc94vAa7xJqTXAlre+pXoVmj2goJ+G2VophGe9ofBULZFulJZxVO3gqKDjUXtV+O6kji5X
n7dkteAcNJP4e2f7ecEfGSYFFDUfwWHgfEvs3vwZsl8MXxw5nNIOQv7bjOl/cOO1Qq9lbL+FU/uk
xRY9U+SMYTEfasZfdRgNJ+jZgrsL5K385wANz9GUPNyh8zu/TUWp9AMeYNPXseHLWdh/j5YeQwZ9
bWUmFstGDwWBdL3QKhHzJmVWYpMlwyoxrBSgWAI9ZGEevhYCbBN6nXo12P0gJefCx0LFwbBRnNxP
MD42QJdygYZA/vkh9BWFwXmEz91SrXlCvqI9B/zz9LSJe5U6R94JeXnMY+F+5jn5pruUK2g1hkII
5Dz17+LiruIpjHuJmH+MTJUYxWH17/gCBu5MjFnZbr1Ia75sXbuUFsrmLQilpIOAk3KfUe2BytMw
tvdH5wTrJMMkDBYE0DB5+4LgN76fqLgaxWKIfe5tUUbrYZuil5/hdrBrKqWLFTVR47dh+rlrKOyo
WNoX0tJYGTTCqFTTqh04u1mhP8QGKLyKiJZj4a6lTKtTV2dAaIVG/2Nza4HS0ZY+sAXFHICesmIx
8SVpbCIxpJ95E4BiO5xgDJZ0nYn6IKA2mGI4rBU+HIu+DiL/g2vYMP01CrNOnS5ngB0wMngxTEbS
NQr6X8zaZgQHGu+zmajy0rpuHzNqS1Nkr9IXrEkShL5srNq+Qj9QcvkOtfRylgEXuzYaNhy+Hg/p
JgRDwru5PoOs3i2PS9VoTwc6F8gurklxxf9MWEAIiC7Nyv2qtzJeEmbALcuJfyo8RAvhlw2FYdYE
vMJGETzayf+eFke4Sc/qk9L8gHAfwTozj5LY/EUN6hSgwjk7kCGdtyIzey746Cdo/ZFuKWmDON5t
n0bfx/WrYH/9kcnWQaiPAU7Tl4H1HlzEzFR1vbE8JtuH8b7X67knZwu43WBO7ny2L7YVWBkWwIn2
WZdPVqdtdlHCYv62GUdbyOjdLJopgymAXkYLT5m8rncKd3nI9HXw+KFtbNwDJKAQHNtcK7D8oeUM
kSnOEryVxdfu2igAANPcC02ajwAiZqdUd5JctG9s6+0KIiQR0j3FsVZaWnFTcLuUY1uQNKsIiP+U
jxvxQmgjFEWTNC53PGpm5vCf40f8FjOswlK7K/Qy1O/xnqTaA6BBtu7CK6Hhf94Cm1cD/my7suJg
LxfMPxBpWDX3WxVcYEUYBTJ6eEuVvPatnwrkss90V9kGDHQsg62Q0qdaLoyHTNyKiTRJ01v/9Jw3
ou6s9qYyBgeq0zwbnpgUrwRfUS06FXsCHu4esv+Usw8OZV+TUcA8hqZmngrOR3NN1SKmYzc2t1ee
7EYSSeARYAcQHIhxwmcg8v3n4YWSsnPO172eRG15ZVcLdeo7Va1VwCL4QUabTdYZa2R+9fr/OjBJ
L5X8OcoZwX0GXH5FWsf35ml8En24tVn0BXsmWtUAt8BL4Vut57vw6BDPuzPbdmgcImA7F02k232d
M2qjpeQ6szjXKbt9a9kUiIlPqQ98TZlqGVkeTchxi3Fyx2bL+mfwEd4ZkOxZwa9SP2krgQPj0ikh
kC6wIX4w9PhOuY85Tk+N4lo6u4FvubbyNgaoKuHsglwCPN1pLWrP0JRflsTsCjKxqqYrZOxjIdc+
f0oqiUKIEcYlJ1/BWKQ7DZgVEfIEIWPBLVYHVfhHdvDUNah4tlAaYWoG/68qe2MbCNXL6pbfd95t
+7cQubd6EUvbN9zkSysSnlMAC5/aNec4ujG0Mi00TOb+Y1JgR+p4WRT00Ut7p0YeYSg9Zsii/Cch
US/JYAkMLUr2WoP8GtJ3YjOD1aEdVXI16/W2iv/mm4HZ5n3kGUL6H0D/73w2NC4584pVwHIpjjLm
vj3BitOTxDMl7q/1R+lrQSROr2wUQbujVoLMp+ICo57OKj7/R82EqYgoUsbbi1Q5020aGwoCMMNv
S/cWXQuQRxeg2J9jGm2wSCwgyxCRG1LZKBdiBVYp32ytQsB024yUBHENKSM2N/sNdn/FbkoIH7o4
cbuKPmDa3lrE9J0B4SdvSQPne/iTgeSywEoH/xa3kuyeLfL90Q/yPvJa+DW2Ens4eMqZXktpJfGp
Vfk7ayA0vei8KQ9zE1ClGpZ3Xs4iDw55jg7Qw7Ot9E5ub2oqg46R5E9hrZZTU9kDjUH2Fp+WvK7m
LSfYDQd+GULCstOexWQoiODzsA8im641gEfse0a5u2rWHd7ugt6Nmsdq1P+9YNa3wD7uFKcYRIK2
0dszH0YlzsjePVcv/1JZGVsm+UaSbjA73+UgneTJ5fy3e08mUhzGAaE0lZxJFPEgKPOqZuPMBTrb
9ct4Z//Jwv+SmkE5ROXCbf0WhJVVAEWmGZjJLYFWPFWJB1H0QXBz66+4lrMq3HMYfnN3a4cIiluk
rqSWdCNH2yYi7zx6Xu5VUwZB16kVvLvM0hWab9AhzYWrJHxPImmzLFxheZ8r+Hrfab/Dzkh+4MmB
+pKScFFvu2UGQuHGAppNbt+NthDF2YMrPrwbzSmofwAFDklABcMF4f6E8ffnftwY9niuezpPAqNd
UnfnW2J29FPNRA/YdNDJaFmqj9Ns6HF4Fnlyrq1QTDiQwdw3wKvvBz5d78EKhfc3vglE/wgeV+6Z
qy/HTyRzlzN1Kq3D05gGhKaLvaSH/XK5VC2t8f7kHlUIjPkCMXmQlxbOjPOsVobY1+RuUc7xSS7Y
DrQPIRuXzhNDqAZgWd0hRMZTfiArkrm9XhjNYauBLy8VnhrBjtSS47B14nGJFwcqVGx09VxjYnFX
LCPF7Ev2eeUvYbWbQVxQ1WEuc4Q4LFBka1NTiYztwuLEv0UefB4NH/JSjavNMsxKd689/GzRCiNY
W5VZNmVbQ96rTgmYbrtfk4yL7s6Yp5ir2Xb7Z0IpYjWK9KdwZZ+oLXrOIpXEQSLX3M+wDfXx64VE
XRlq6SCtS+ugBCJTyFBmZHAeJh18f1EFMAL3/EF/UK2dbacvM+daBrFoiN69FE3QISGD8TikkW5N
Tl1Hd4Grff5KsMkzkQ6CXa0buwhSh1L9J/II1OTPbQvWehSSmmNebz4/AJIIPjL+BT/EVoYhz+LH
Qn3PKnV+nNHU3a7k6dgzKrp0JtVZbZB3RAApfFpQ/AdJqhk5iqASVsVNtZhZavuJd9UF6BP2gtus
dCDxW8Xozf8otaasHEMZKmxJNA7ZzxbTiGCJQSDkjVGUDX9x1KsW81E80OBjdfX1OIdXW+7WhHci
dgxawxuVUpKBL3gU9e666+//wrwCXRxYZPPqhWSWKlSvCk0YKy5A16kmjPfFqAmGvvSg3+tDSJEa
15fbtzR85YTRQ2Oa7ZEfVk96T84SMe0cyEvFiaQs0Z/MTJBv9MP6vwhxN3zGyFaUJ05TNv3YR01K
klgk/4MAlXc97PWuGjPl279g2XOndrDO80JfFKnHq6u+kQjfCIva2kJpaqoJRGbwhs/24fkuY8k2
menvGJuV+pMuQSKtsrDRLsaDUAAZUvXRlCgW9cy0Tmj+3VoQOomZTc/XvL7EXp+q4mGIGwuNQvwE
jW8oU7bNhkt3Hp9ULtpULnYxX2j8e0qUNwXeYaQpNHjBScyA56uG51OtgMlrFEBKGuVuPObCHyL7
yB9mX8E6awqdinIhU8PHVAcfwd8GO/hAaE5rgVAhKMGBriCiCthTqBIC4+/ksFTOvKvuCd7K0Zdi
oz1CV1edyyuRNC8s0njOVtk4NUxJZC8QN6Hx21x78+z0xxljRr0h2fSSmdLjWgJT1cnZmHUomp5I
zBzE/xIExvb2SPL/I2WYF21t33w9f0CnZtilQM7cHWUxZ0CVh6Bb7XDoy5Yxoeuzsqj2GtcfjAeF
8GSPO1BHx323F3sFQdv11M6jrA2KaYYGPtXDPoSL6oGEid0mXpIXM0uqCiNFy2sjXmhMBO+e3zR9
p2kRQoR4ocU6fTCcJE0q+CUZJsGX8E4940u286CmqXOv/gEa8m4redB8ZbojHksDoVEI4jUw5N3S
3J1NIb4uK0OfPklhRvCuQ3/Q4G1w19NYVOvVTh6aNC4/8hj+2cqTRUHe3i7raHXLcGIJkwUV+YPU
+IbXsG/B8jD/BonYj1eUDztZjoVqFr70zHuQ+ssDKiGiupfkI56eFcKkxwuyXp9Ci+6hXbYfH7XB
mNtA8LK4bzfAC0IVlg6oI1X/SIbV1oZ1MoUS4PAOKGtcw0sr1grrTSDUStMyt+STcBtwsmISe9zE
axYGx2nZNaX2xAwCnwdN7ZDBMBwCxs5no26tNd9HHTeulnRU/Pa2r53N2wV9ZCTKLzAbUjn3owN1
lkBs81lzJBtCvW2R3uOLsm3HqiIrP30QxTGa+DYerbYo6DLOVBOChXgI4y7iSbm+kSKEyHJZnvlo
J72LmfLy6hu1rCZCVpKqHV38YOVusesPyXk2d+NaR8sxITwMo4Hx1zSctCFlwXKlbjhAn1W4vREi
6ECdGLFn/Eo77hu7kdmTN3lFWyzkYhuAxOJWxb32Z5G4X9BxPH//EUQsXIb28AKd/TLtNJ8RwbCW
y8uT1I2YNaTj/10BZv1MMdON2Hl0JPXaHWEROtM6hkIWFl7/LppdJ0ekjqMA/PU0eRgLWTl74Y9j
hP1qqogRUVgM72ESjXgmQhuE42Lh9rb/Yrf0Tw1mi7qA0DEcdmXXi+Gm1moeceqzCiLiZbaxuRT+
qsu1psDeFAzteBUonVFfHxV0+x2z5RTnTfsLld3IdqkAPYnhXSu1X5a2/iq90Ud8bkGdaaPnE4KA
+udE+wn+YgtoQxYk0ZiDARdngzB8MBlm1y1A4/UdNL5YSI86UArfCVi7xh8jFA2/x0W+nCuFqxeC
mHe7KtEO4jGuavWNu4P8rPyq7MVQMHx9UDM/ySGIqoiv+13GyE3AL8awpH9r+qW5cZMqTLgBNRU3
qxYOe3LmzJoCnS7KYEdcktptT5dA6HCqZdr6iItf4O2Qtw1b7Euwp4v3UAp7Aulmth9ee50Lqa8t
Er783gz4Q8+UxLW2IAkKvHJkIiHpVJPn+McgG4g9m3AWI10xmf0m8sgwCrLp54Y3OmC43amzDQ90
Ps6ssaiJYEsRHidbTcp/1FQQd8g93o2sXdQ+8WWNd8nJpy9KaTI0gHApnrjAkaqpRjPshOz5I3tq
VI2KmDS5hCXWy6Pa7PAm3uRIg6Bn+u7wOLvjW28cB2uoyhwDb/e6nDIMAG3G2/iapBurXr6rCs+6
oPFprG950TwkvmnCpUA7aWF73GWaZd68nLB7Ci38tnYAv0X8iSlal0pLnfbxZbv2FkAA8UBcYXnc
ke4ym2y4l5N/vNvrzLHGLYNARVlOkoySxL6JZpcQxma2Gevo4THB2go7LerUNAPcTZQ6c8mSYqJO
1oW4iAYpx3yByttjKbhGybGy+mhtSrrPhZdb2/q7A6VoO/U9//XL/hDm85LWjglUTzRc5ivNtTpj
IdU0nLQpbsUVP6fviyDujCJsCPjYp+PaAVdD/bSV+cYwLNrWCKlndcKgDYCY9Pbw79acT8ibu+iE
IAsENjKc2kquCeCppOZSTAZFhOCVQZLHGJzkqYyL/LLG/PmenkV+BOOjHWZm5l50GMiuisEKNqGR
mkFtEUIzagxCtI2Uxh1uO4Uolmv49wsZn1KzaMsoYS5Ty4L/GPYR+nUeXtuc3fMaMcIao9w4xAVW
2FuHkmuKXyH4bIWPiwE2qcNd96x99/qldR4iBTP561t9GHV3nxDVJuPMDLq5w6iiqQ5ATZTiypWr
Ikkc+vQUDHXA3bBDyVNv4mtAmTjwnbYrVDNTU3jSPXMf0Z1Hr0U1xDbfNiQfWGkjfCb6qlnitA/r
rdsxx1wC0AttzD9qZe/pEokiNKEzbUOyuu+jQlNO1nvCt1Jth/mazlIC3hU9S3oQm2MObLq8rMyQ
Sgdmt2hDjLNubF+PhIQEYFnsaiDD2K/OftzqF2NACXqPHsGKAiNIcsIYzOstd2TACDIChFZV371F
hn8WxjzC+C6ED4DA84VtJfwaw7GqqpBQ59B2d7snG1V5DnJhXfoWecNKbbf3+e4hX0FwSXOMjLuG
MsQR+TTxxytsY2RSfHLkzJA47UtdYTt0yWtqU9xbyEi3cR9f/I74dl4FKa5+DnAA4Gca7XOxJx75
zgwybWB3pMRt8LWOnYf0pp3+4dstd3CLQXq+A+e1/gvFiguohwKAFskYV/y9inGt2Sb6VMbpTRIO
0sPQAMM4Kf71rh9phpdDBQ1qMC8a+9umUuHgsAd3RQCMzB/0wWt/COGOHCLspNZN1rLRZqL3o/da
lcTRWIZ9ka9KtTv4nkjaW5BHmsWgkpBrrui4SEqAsm2bAA9Q6XSij5T3BwPsSWbW+yxN+sLPmuqy
a6TxN/4P6wQKKGnZ8BY5eiY2t8C5S2ZLB2xFBeNAOONGMBpYOLwvKIlgifvs7rmoD+VXdjg5bfrw
jX0wkuL3AO0iC8EneS8lZyEVIethU4+GyoceiFL38b1Xa/caCk48Tku7IqOkF08IsHO0K2ADtxYA
o6IGJe8OVg/bBhtLosYRq9GnuPqmsqNJTwKZHp/i1Vb7zgQI96s7EDmUOiGPtuvtY8laPUkwzWbz
piNR/A5AvsPw8yBhLnt2s2WPWc8elAEKiuLlk3ywG7G4+EjPZMiK+jCuDhw6C1qZJ9Kb0WTdJjyZ
F4iC3xR7vkIg9DEeOSq+YTWP+vdIKyvAuM3ofYLJJN8Q2C69xQoS+qqxaI4KQQ1IhewkTY9L8sTA
S9Ypji0fvQJh3gGQF9f3NFkdmT/s07mGSd/ftktqOLZelSkO13w89MrdwRozXXufSooHSmVo3WoL
5ZetBcHcHPBoNXFNHEzoeZSmqlOmaxFFPyTCCBAN5TOKhbSzPBaOsMANOjT+s1AMWXOmDHzFKzNR
HZStdGwjAh7ekuWYxaW0p+OSlfEPJ+hJu0xBcmux15b68K3Kg4FGOgfhOKHzCDAIeefcxiXMcbUE
fJjOayaOkcituFzJcnqF7MoGRfiDnpg2IjL+fbk3C/XQo5JAIDpuFufHCQBtjLCXXVFRMMza/FRL
c8dQoO7791mWgNzrZ8JMwB6pUQfhxxtly0yBtHHM2/1PdVWHxZXJKWBq9dfUK2zRVug/VSdrMyyM
Hay2e2nCPhq1d1Qkeny5K62ckKA7Lh9/BuLc3Di5WQw/ZMipP0D3iEu8voSSdtree/492QZovtYF
O+nL2pe7D2tOUUOKwYazQtPuvlp2036aDZq9jQDfg4beIFr8+Qhy/t0dlD0YfgeacZvCL3H7j23S
6bjc6Q8pHkIyd3JMbFltYHGx/Tm4KvpwyYrJ4Ttn7gpDFq8E1yd+kmtexQbrJ95/HTVHFvDIeKx9
agU0UHvjHS92z4hN2iQM70E/rw+Rkmy2Za1tuysp0mYLjkuqz3Ht/EeyJxtnzUwmATJ/ek7yoH5w
rspmHRA24bEbgsHEl5xpuh4B6yD0FOywj1MtiyvaZ4NBRZpwF2En+SYQZz1z/kQSznR3vrDw3nqG
6hIVCVwwmWwISuBoFDwDp7i1xiwRwHmeEFM3tyr38Djjf5y4phcYSlhWEHbFkVblXxIDOA0J+4TT
IHBZh9s++wvzbklvbSpg8UC834bLsB0kF62tSUEnOwXZdOb5eOO++3T+DcspAIPy6QNOS3rM76l/
lLvozGqOYz0nevBqyqNM9koLsGLMX7taX9aai0FMaaq06/JhG5t9WuyFZt8hwK95SRVjcL6YguAh
oVTHh9QE4L9TzrylmR7uRrzNqbcXfK4eWUqfifS23mEN4RZ/hTHMLJCv/aTTPAshdHBC2P3BPqaL
CRRpE5GRCAWi033PgcPM+rL4tENtTnj73kYEOuyjHaYC0g5slvz12GjULDlHgjxqk7ViUgVetxVn
MNlYnW7F/1bpR73Hk8ZyWadMRbeUoN6AEQm2jjbIib+12VEPeHojpBJeMprCSgiDvErQINjHax2/
Zncac33xKPy2YQ2U+Kf6H5z44Nhu9GZDqHStoqmMdotMPGScYsHV/39mTE2AQQWXJWSRXM4TgUC8
ttuasJq5eCBUCzksAxXTDXOiAsU7XIs2Bg8xVm4IR5k5U6eWlb5eJLUPS7ED5kK1RZuANBqBPVs5
S2p608SLi1w9XUtfZXuoIcXiC37/DInXxVdf3hjqH98DtvekTX2o78ly+9B5ucv6xEb58Zxnpuzk
QYz7B45LbfpNxfbwhFXNtMehHxcTkWh/5qDeRAmdVrDdTBxOkJaRVPyH/4zTgBAsvBxA/lLpsfrf
/fS9TtjLh3+tqK7NlesiMvJ4l4USAFbIyetY5OaJO6Oz5VQ8trRL0rYEsQ8Iia6qOu+pxdPbl7Wj
94ccXx9xMPkgpovV1WjUHBsIx6FBNTUQE4CCXcFWxCyRYmBZm64G+KBEbnlpXrgFsgvFo/ScbhfZ
APfL+46TMJ3vxMOU3k3XUiX+b+TVrC/w8XUKOAMCecp9gC5BIo8OTn6MNO046QicXCGkmlx7I33Y
X0Wgw7HlEh+UINwTqU6J6UewaKEd/kLDZzSU12SafcQnHfEK0k7aiAljO3BPhTgBVQEexgL+mNY6
+kI3uU3CiryTTTT7yNB0j6FrpX8sVCtjOaqYtL04ynN2fqTZVBZHbVkKs9UJLrfi0sE186xj42sa
h8YYWxCstds0e4MmhCSumb2O0fguNOQ2c05dh34qI39xdCrm48kpv0famFcV8i2tHBUPiUOL+Qg+
iXJ9RKfrVTlpS/APlhIjt0YX5b8xGPexcgIEe+czJ8Z5TWdo2VtiFRvcx8aWEe7TM4zKvRXdrd3b
B3hEu7tks/fbwSvfzr3sKl70YKqBiB08QytYXYR4M50nj3j0mmGc47OUZAUX8M91h0s+P7/joY98
L/dZzJ6s8Q1hM+9Olz2oerDRUZfL2wG0fcjkH3n30VEwj91kp46C1Vdcp3Isv2e7mMd1FfP1sj1K
DfNvjDRVIfB0ShM4NyUu+45Q/MVDgUpeXm1ADP09AgW840kYtFg+jRVQVWJCy1EVcaigfPbYTMLK
1XZiJW2H6FNAyaLHluw+f9hf007m+pcYdC6DImAmkPmPyx+U8CaafnF+fDa+i/rVcl/3QzG1J+8e
5CXf/ag1siwZMRPnEVpk4JNMmM/WfivO2EWVqc2fBPIbYl4M0Jv06MdsOmo42Wvc8i9zTsbDS1gV
zSo7VrNm0b4JPA7Uifwzn1narop7nMSkJU67XHHhbmjOVk5PFSwkevS5LgA6bxJk5uwR2/awgRRn
EDVs9X6PXLcZGLgDvvWaA3vFWX/969LkDpla77cH+HIGNf2qP3FBMjdN/N6qnsaWNsRIesX4dhX9
TUr5L64LxKngRM5C6U91kyEA4FqD5RWMrqKEC2nKSzPPDVBv6B5mQTYFxIkn+LIfPxSQNtqL83FI
KHgL3uwjgSbJ88c+dOy5ndLoLiUo3e7o08tEG9fc4X6V2oMifqBLQuDHewbOXw3ht/VdjMMaTEDO
osznPiIyZBKYleTQQzJgyMRQuKAOMldSDuIKH8obGQIgoGfmkuc56znr2DnNh8/dGE4rhJx8GbJX
xrY8A44XD8vNCBhHwqGrNPOY/KV+QjMOgoxd66LeCHu36ZXNCvjICwzZzBlHp+RCuzHMTcGdx8bA
F1JPd0Rs3mnW/XBRytuo1rhisl45Ocl102paNS38hJfUTA5vygozvmqQUHxrtjWf9m5OHXmTUM4X
SI4mtHu3+A1bSn1K1XFfZ4YTkKKOuHAcbwwXQqHbU593Oc438Be49op7BGoL7gKux9CKDCrknqK5
dQjLcTpAp2g/iZis6bmHjyunO0H7hCnlGp8cq8UvXRITC6I8wzKTXWT8x3KkueEvM3DJEtCfYjJG
KeZcZyxvPLQq3ku80I3bJoQzjKtasPvMpFtckfj5XbIrsuUi3YGja70E5JX8Eh9Iv+uEtY7eeHGY
z1UUNWcJ932cwQAa94iabRuHk0RzlLfrcetcdpnowQRD2C88/Xcc3AEgnSbKe4iH2alAyxk373pG
8y8ge/vdAGEml7/SS95IE7cHURKEazKtgkFg4oYkESf0OrodRuVEPiVIRB377t9cxIxE7ZP5RCQV
ZbxwMWFPMWEwkBhDaCaB8AzE4EeIBmSF6nlxc+kv1TfGyuwkqGiijJgSkGWZVgmVxBFe/8kjWuY+
xsCakO7ddsZbmsiifPAzNDPIJQn4fZ4tL6CfCfw3RujJYMX6W4otarje9BoV1yjo91WxcjFy5OWG
JZrLTUVVjcINeYDBnDw2YNtN/22QvDaKRp+CM+ymZZ5uRSJHmqH+DIZavhkVWof1xjoiKalmMybE
jIwDn4NVDBTTa8FLBVKo3mZ3eWptKtv7IjecigGTU/1OScEJVcZJiiJu8eIPOFrVSg+WjA5wickV
czOx5GURDrVlmiq0ICcp5rAVMQyPD9EwWJjhMfPzXZhjRnDu2oKer48iaGiE0ecMYWVFgiWnhiDj
5PCf9fC8/4nL5PqwfMS9LBjuIS4Yk+5keScOM698oBbpdjcTYDl+PVMN+zxS8eKDemdV6EKhi79i
XPigVHU72BM9XbdYWz9rM8YMQCJ60Vq18zaoglJ949rJPjBvju6TndwPhJFDZToFjLg4Q59T0dMn
wkkl0wp2HqlPMR06Y5p7k8kclT8yisqx5tJwgJIh8ClaUIZOV47B6eWsaoW2S/kr+nhl2WtOJuIk
G9HIe+ZiDvAQUb8LNrNS9SKn4Hv+Gb46g5+j2jGWwSjxGwRN35eBfHGRANTFskwVX/qtJCz3zwXo
ciQRQ6wPuL7gpfIkcZQ4sg68llUmG8iEj8D4JnJiwjrd8BXCTMDT7LC29A57534fQPt6bDCzdRee
64H5bWgv1ykUFdPC9JBTe+U/0myuRWl0R2V+sP63y34UZOV+rHH1z5xqQBgFtxpahthBatUt5O3q
yKBr5Ne8z1/gBlZImCPq55krLioKKUM9Guej4aFG8u9QvTZzz9zxni2WspSD/RXJpiMC1wowijSJ
rp2jh1q9vPmFyBWOJXDZcfN+3fLCHCdy07ECeIvjVsAz0XScvss4NGEIHURVRb+k7FDU77Lch1Qj
MNyqeLL5n3XRgkVBx3bmjpAQYnm6CtZ7nviJRHUAFipaj27dRvH0SbR8R38AZYTcjE8ExJgUV9OY
H6ZpYwdXZYC1dLMdpbw7BRurGvuKLbN7eV/ZjVdwZncAIh7HCveyeZTTVhzsy0ZwJ+JqpMY07ceR
+1+umaCD2w/u5Tl53KIJaI0zHUCmAobWRZ4GPcUs67pjxnmfme749oC7DF0U8C0NBSjPKhhw2RIG
Vt1LlCk3b2FS2Iwhexzhxcs4pNpJUUuAIwyRnXH+Z+XV5hZD4aktg7a3jHTi0Pu+wpkPQiMG88JS
VNZNBeH/72lo2pz9EPdMMSt1sDK1hqvNe8Es8Jp7zaJ55Fzi9G+4IpxGSYumdavQsLKQP7YHZqAg
mDDmd+/nPrFtaFRk+KSy8qtbCdMWL7csFc2O2inlMmI0ZKHvbB2AEs6bxpu9Y/5ljH0Ogw7PCS/+
uKbvgEmBzc8UT+Ci9HWAnM6lySpt95UKlHzQfy6uopVlGODujsl9QgDChBPiqT7Kbv7hkhmhTxTC
7VKw2yNYZnO0VjlP1H9i29Oxs61hmAnninUQjO+EHmGTFlCqKGunRzJuyWBZmQTtjhmPCnUZNF4P
eMrvzx1R9wUnKo3sASViSoCTCg/yYQxoawGUyOptW6FOdpp9gvTuQAxTQFrdX4SqktP/QhOhPWPE
joQZ/2VkEjPBqEKuqWZBNb1ivL0hVpWkaoCprNlnvhC/JwVMqoJaQUx5uN5ZlZKTuPvkAYexIQok
9Kh4C+wqsiGUXvzCwQ8TSH1yypSc8sF8aKzjJjaZf3KPq5ygXCF8GR+0rZaV1W0lp8rb+DrDrdSL
1DKBxy9x8vPhU9SihE4bkF5nB7SyXXlNp3ivp0D4sxMoGh9jg+xIhZifkeOQHEbmqdKpn6FtmkEc
QFwffi+wsv20trM0ihiNCdW2rrwL7yT3oCfKfEVbQIU5JiQbbbf0cbQLNB1mY6c/ASevvKOl1KgH
yB/ZIkapXUK/SYKZgOuBWG5nSpstueyEv/oGXwMDfAncuZJxJeWE4g1pTiI3aN3pPXdrTt/UysH8
kstepWB2svPtiBIW9VfFRtDlv4FO1JQf4MvtsM6h5XajUBUm9nYrWWTbiHDbWKqObEMAsfO20vKP
omtRCWylxi33em4YYBeo3ms1uNYiYOiRCpko8tiySNIUZ6Q445PdWgdOyiFYW/d+4q4AR/ARFI30
/UdaPdPzLb/PMe8wXESmpX73Y0OZj2zy0TqDtWd87TaMKZIhdwfwKED4GYUmkx2Pn9/KugMQTOUh
W+5ypJw4Rx1zZ0U0xrZGNf3M1795kuwha/V8J13eSwXXIXZMDrPNiQeow32Z6D1ZnQWBKp9/a07y
5V3UZnuJ+O4v0F7EQliRMIKLhgrqPRl/ZKlYrWPqQycy7ZFUtAi/igmyC2JkuFPw4iDffx7uuwMX
FVDFSNk+1YRXhhfuq0akQ6oh/U9AZh0VRYUbxHysWko+fZkeBinuQnZBoLFYmYEoepL5SB+/N3EM
dde7dn7ju8mse4Q8ywZSra7jsYzEQKGQP83/RXBR1joFkwn1Rw/bOJ6mD90ZNbhAevVoVXiVwbip
k5W3eybfZomIDweAob0XFy+15nmv8XZHBs5Q1+4MGtWpK8q6hM/SL0vSRl0sJEqWGuFQSp+WF9+f
7FJS5he7LZ1UrTdxESeMeQdOOdV9LQgdZi8jOP1XauGRytib1nqTJEAsf7/ylV4LFhx9kRvB2Sbp
KvjZsMgsGKbWvpIledEJL6GaBUidfo1rQlUcRZHOlPtZ+wAuLnHPH6KUWxwAr7iMMGFpXV/stLV2
1O9ZmYhIHUvv5no6JKmlvVd57xDTur4ITCWyrzOLIIjMW+G4qJzAzHSGIvXAohd0vT1dKCUun9pF
eUxuJZKVEe9mtVMltZZsjgPUyyL0rERtmvjh/F73xejWYb0oyOaclFrJBeVbc/PlQacA5B36Gemb
lNwFyBrX6pKKYOuQBVqiZF6foTR7CQQJ3YHOu4xkVtGi4iROmnUzrVNvUky8QBqqlnUyDBh09JQ/
8Vpx4296LwcUK6xF2Io/dzRBjyLM8gnmgzOrAF3mhoSFfBOMWQU5vWDKIvcshFO+++NSBi9tU6aN
ib/pWLzBLCEcAooH9sWasMND9QURJ+YOTPK3UPc+I7852K4SS2cCnLcTc8AfJOO9x5bS8yshY8lP
+eDNPYZiJcJf5Ze6doEq6fg1CfboBUei3yjIVJmgHUkf8yb1JrEXCWXgosbsCD+EDZYFREcifpgw
3EFed7wrJ31ueB63kAmqOhM6iMZrE7/DNVwvH0U7qEpdWummw6uRsWLvRva8znoLoxWdkkdmrlQ8
SONkhgUcp5rZh3zVflxL0N+8qrIt/Y0EesjjV0VUIHpWW09UFB532Pqlxu0e/7JoUgX3Aw7Gx6JP
miwuQ+qpuFLiFBdmIkFX7uuRHpbb3zVKTJeVUPGtGD07v8cs19+d2EwUb6yNII2sU9+K+gmaxHwy
Wg5KHs7TmFSgs+sD+Db8dxotfOg6brKcUB4+ROVuXNVxIHNg2v8bH7CXqdtogtYjaX1YIdaYEJXp
2K5PEWMPEwqmse4ofH7tj8d9MRa60oS7NCs2MuWfeI2cU+w0md9K8peIjLYcDwQml0R7UHS0JX1o
IpyMlIHXKIrduNIFwQ7iwoLQilNNvm/NJ0EMfyyfwSU7g341NTEZOj3lBKNDbcQuejK2nrOVWipF
L1KDmknRvWgBUSe8ZtcUwYB1YPajODAM8ePQ0fEe5u3E26/DrOrwT77pS6JBnWrHM11KFKRuRrJC
1Gwq7N0/dExKrj8etM7BcrfoUMr7CX7Qph+/imz309Qg33DPJ/ttgs8iue1+oEakuzDecCrMNFHJ
3V4BffSPELZ+gsWH7ljGFcpAOGF2WOeYxtJU7TN/X1iOKXnUno6a5Txfxq0us5I8q1Ce+gTPBFJe
niOpPMHUVRPZJxPrbOywHPzx+r57vkiMfS4xp5TJeGL2OHomWS75Umh3Iv2z1Z2eCMnLZyDGT96D
V2AwVrDiiO47skdDU2+ZEdJOJpMTIAfnpQDzclMEZJmX8rrgiBJ5PRL+Nw3ZreBymWT+Uyejp6nc
RG7rbBdIbpoP7GXnF/5ARDbAo9LcGpXtICCVr1CwI8OCAq5CBENc2BVWGjUh2gromydqbBWjNXHr
W4fDLJ7+D8Emcin/exZ1dfzZlLEZFMavEgIE9V9OczmszIDGI9uDddkSMLyKxeoGmw4TI8UBqidQ
Cwqgw7MgwaCI2cgzd/z7oqAS3MXjQxIyvFgTC9QncI7d8iw2n6a6F/GU3OvLpcogLqQ8sm/k+iQq
7SuHwl6CkRSqVVLP7YJhoZa3JpCanw9yda8BdPX4y9EZRpKh42oL3QJaobqN1tdEVttUvFF10VIu
jzdX1jSXOZMoNnv2rqfL1KSRQHuIKdqU5dyjS8w5ztDTTrkkPu3ReiMwtafvq3AoWSZecZeQF9ky
u/T+v240ezAjbmQm+FwoJNj4095IEd3E9Rodajvb7rAw3uKQNt1PCnoHePvq5wNVLFaJUW//VWOe
Q5fts0SZH43t9wfAQQDWw/oo7g2JMTltEqYRCojWvb9WglscpYInP07r6iXWRdw4JZkFgwq+PO/k
DbQDFg45YCuhCIjV1YzvEaiImzd4rNqWLzmcTz+02OiqpWxiZLoonKNul7VF5q072Pt2QP9LYi4/
CvudNMIknz7XNNU6ct7eCAmMpYy6Q94GF6VfozY7xe2Naq3CMV5SFcoHmEKaqrLjyMQ5B8d7vCgF
/qycu++fICwMKtbgF2KAx48LCiHaLtAS9bFn9bDaQbLG5fO6esxaMzAvBqzDKFmMuxPwl9OO0MOZ
d5pXYu23heWVgfs8I3g/0eEjPWn7ThPwjjKw2vU4rEqUIOIpck6y++zBX3LXDv2liRvMvViiQ+mn
V34qAxZ0jZAcUL5HOVz+l0AWQMyt5wlqbZvaYc39U+RHh3zLRk/dB+qhAeGr51oKJolv6TDpaGzf
AwxsM/sxopc48Acewpn/eKrWDnmf5YdB8XYIcdfW1Gbknzm77BxOon84w3B/Sta4JDsg/QEoQEXu
ak2teZvRhou4r84oGr7e/+DrXA0pZmfzOtVXWX0JDHU7lSSeR9U321XUY7IE7t7c/BYXPDdW/e1F
3If9JpsRj+yHsC0rMVbLMzLZQ28H5DtS4SDk0Hti4VTObESRpw7B4RuzQ/JGwFi3eqIRKEvNJQCz
gZ+QAHAEaiukPFXnTiFg2enNMkIlDRYxRveojYFeNyfHKZliFqZ1M1SnLRvhZCs+Zo+8OyyLg6vd
KeAo98m8FCCP1+9fSXLKaz6/OWUv5ZXJITOojWuKnSGELwDsn1y2YmeJrH76Db5NUy2ZHXVPjBmD
LD7agrWcgQlfxG3k1pWt20drTIR8L2od33XfBw/zf26d8Fr4Xnjcq0CbESqkzyYvAKSX3heHb109
mE6qRVB8qlR7XiFbjg6VtawtXluv23RRYxxdctQDM+bAID0aMqQe0j8LsutYgxoMEZ3YFAFsDpiW
RkkTot8WMdq0AO/GTkY+95HSp4XqE/5hRSGiiiL4jlXLPzlbDsahV3LNaEhv+Gh15ypppuQXrW7h
/Q5dxu/Z8H5rvUHdxMqjck0gFDghf2GXQ2zCOXOjI7bzmLgS0DbOyXofxkT/jpTIQTqD0N3zqhJy
2FYt0GJlh+LWEOJonuZhnofiZKyJGueT3VQCrR/LyyaHQKSaIDPrYnCxihiOJ4QyExal5uo0NVi1
LxJ9HsXdk5TgrVq4Lm1fBKz+I9ocwfrex7JXt9XSI76rsoVLDWi4zLAe3tr80U7p1QIX0+Ajo0cB
qlyz/K2/X/ks4LZWU8zl+v+V5mAolNaUZlnmGUu9VEoG28U3cmBVhLIDsvUARUv1++frvhcrnDyT
/wuTXfskVs83H4YL33p6zendk76DcEdnuvhzroGIOIJoPesocvCA1VFn1R0xIbt08JEp4ZnRBa/V
cVfGxleZnbToQI5zwNsr5iKtjnl1eKu+q9/Hi8oG4X8ABJkQ3NZlQIKzSfmDfeWrxRUzn5rbTndh
q2vW8IRdFXbRIwAbH0nJK8uKuB7YJgijKnNOB9q8kf5M2CVU/srk1dRPLANRQZvH47ErCIh2183h
CdRGkhtY8/98jbe+f9ClQM1WPdljPv60k+1FhLbMnTe1o/UQOQsMm6TxEKZEOK9RTY29KJj8KBpo
RYbaUw/f+JMFCT6BujuVN6IPtOpmPlk00HZb+X35oFRRS7r136TigH+LC8/D1MtWRLuRos8WInxv
xuwHAzFnDHrd+HuV5k7lMLLfOkrUYlZG7m99pSnf6mV6elTaPdgD4t1g8L100htQtd4QwdOOVgri
WSTySkCiai45pBdI+CEbSFTvpq48v93DFQBWfuekL9lCcim2yBx27lIEWAT8/sXBumOGTsuRvB8d
7O0oFqdZURcMp6BQA5nMgkV9J9mVqljt9QhCtbgCx++6qg/nOn/J/aG2pPL3IHN8S/r+QUfaUbTb
ZiFLow9/d2ohQFdH8lypSaPkOszRTzvmgKlMlXv6HEMABonUjYANIsBRzeui+ATj3EFzLLcF7sdz
vYe5tOL75QrEY23eguBNdMvbmd/9fekXbB6W8gxT/2p+LuzFUfFV/cwKfhXRwfaLfrdHagsqYuk1
Jm+70OQc5bffIlqjONldF6bDwH4ShLxdQ9kDKnNdBEb4K3O4BvK0PIIhNc5H9qwRJVxUFRr5FGIF
BzDAgDKyPRuLuYwLZMb2wnd2NvnzrpOx9Mzp/6a3+47dxy8wO6WoIcqraTsch11EzMyyQtLmzmuL
7iR3unfsr6wdevs8GRYx6F+beWHNys7erKmX0l4T63M56P8JhVpWzTYyqQcanvHNuj9Zg22UlQCS
9QVnENTrzyx7XeohL2NeE3aahvBOe2MmmhB6RUivgPaYE/ZCvlXG/358kNHeujYxFfJixI4IXHU5
EojWs27mJ0pLP4HirGiaeE6JiGPJ0t/8vHm4SdQzmzqbZ0Hax1ETQrTSAP3jgOvUEvKfUPCOAEYr
cdZVgVEvRtXThOM+gcEDfmW8gTspuDHUm7spezeFZj3N4Otomkj9yEdvpRcqWzJGn+E8SLAyT8dE
GzBRNWMPe+XZx1NYHcJMi4ZYiqImJspSTzYTIQPaARYFplJV/miD960Rvx04J3ws8PRRSi52wxSW
yT69fvhJAathcbVB83sjLb5i0LZQVIgJ5PiqtPumN7PsxqPEl7ztOHi1KODyDsZ1exLPZQ0KerSF
Nwj1qiTAvIi7dabPRu7IYt4ap4wJhfEOG/AQWtivvjNslVrQtS+Boy+l9f1GPk6HaRE9A7qddbTI
ClLSxlXtECtcc2HVNESP6IcyiqwfI/S60ndBjOmbp6b5AGsCc3hCW0H+RDGIuZqcsqCfc4dxLc1p
3GDr3fvghe56mEcCohoOio6XNInAHWUEPKlp+Edth1+FIllPD+7+bPw0Hmaha20tk1Vlcz05zLL3
UVaKGYG09IqqvyMsyFrAQlKZexe9c9I2MDFemSUJP9HFokeyTURZ0fYc+RvX6BwPUns57eXyHYS8
Oa0U/8lzMkSJ6nlEujGLdC5mAJjyvN2jmQpCiDWJReNlhwbk2b7Ujr6zGs0dtkib1aaquDWvGCdw
T59YfRdbh5DBmBza66XVy3d1lrHDOvhHx9AYA8lXOd+vQSBqS22rR0xhuMPa5cs8zl61PgHK6Wqt
uMpiJq89+VyyB7nbF1hoLqZ2WLo1h7qtWXpKUb2m1Hywsq4hya5VnPWg0Bap/2Ct4hzk7ndWget+
2Vkyh9qVz0bzhswxIaJEnbz0J1Ihe7XiLrfhWT0n/3cRKPdp/q5LMLPFPH6TIq/jGzdy709xd9pV
R/rh5cv2N9Oo5MaMufwqkvfeY0mh9nEivoFPUV5nnWINLcAgGzrgwAdImPUOjf93vg0O0ho5u4Ca
6IsSxN7oOBWX51GwBWhG/T8XYpPsYcw8y3e+35K8nSDqC8n7/axfJsue9nAUNUyAJQAaWLyj9qDV
fU5NlOPvEdFSdbG6Z5qXx4FBs49RCL9naISQ+ddVfSsV4Kvn5UGZP8BUlYF5pgWh+a+/+j8SkPUX
iJlRLOcrgvIxOhKGmrYJtE1dc/NEWV8vwXHjbkGmSwHX6RvqGLRUUXhPGCyuzDlRwyZvrloLsDGJ
tV3H88rMckiwQK1Oww10YDKWJpHizmSqLC/Utrz/TXgRGRp0r2qA1q0HC6SUmztVogtZn4G3zSvO
9O5ni+K4qMfC/ofgiPNpA4eXGRji/5XdJVg4kYrVgVR1BzZxB9QLG8LJPs8ISXAuv8z7bIu4LRHY
Q3A32XNEY3sm0HTH/0HTQyMpitwAdwUYtdp6L0HffMshb8/vBh9WzPxRpnA8cpQcwHlWJetr8rc2
JFM4uQjqMYJuhkMg5QOBec6ccz8DYaotGkU2aAp/3Ck3X/uK+Z0gAkSPhlgjyjKFP9uKQPScVwHG
tn9j4JpDnGFy8f9+muhPNYq3rjPzvQ3arrbe8CZodJCYQj1LD1DPpjbkkhThd/sjOCwUdFVhPo5g
mv9DmVgSLoLy+qqjdb5qIiVpdEC9Yp/s0EF82SVMlhnq80EKh4XkANGmKYovgUGlyCmedbKTFnI8
209G5xTskFIwE6P4W5lGX8CLs3gpo/6SxvSjSzq2gb8CJeJfNRqVJnjETzCA8sr/dTUBWP+609qn
oxrYYArQP9jYalftSIs+/NdjBjL4u42MV7rHTSjeIum585+B5V94uFWRx+XGjKAE2AA1mInFk9NU
/srTnSrFUuRxzGmzPgwV6j0SFQQgGjzw/uHFakT4o/POsCaMko4CsZaLw2uQneDBQhkdG8dV/8Aa
a/YRg8uuaUOUgLFLmaF8QWbSOWcE4HE18MMFm/aVpF0CiiqkaMnLrK07bFeqTJcZf8Hoe4VNc7nE
VQvHJHu3QltA9NWnnGZ0kZjLIGpVfBJUaMuXTeggZ9abI5cNglqn+tJIoT4nxUv33BUWWSBBUBMQ
ZKWQU9zmV02lrL9tTjsbOlTA1bZ3LV4tJbt0/RaHibciKKGDPXp+Qgjzw10Oo8WYv82CiLp4mK6O
wOKiuvSeaC1zUbwHJ/rI5ILEK7q5x2zS8JPMUxylA8sV9ejr4wEGsc7PpJ/1JRJ15crkL1O982uO
993tsk1yOJvK++fhrArtaJebXs9WJ0P3MQCMzSJRPeKI2l1o1Xt1qjiYPns9aPwc57q15jwzycXC
RpXf4bPisaLkgnOdrP67+ToPGuHV9J6Ry/snYvj9lSNpWpT042Ij703HazXBEVSU8SzrlS7MVm78
i2Ccm016/t+otaxXxZ+zEEYWE/31VcbJo8waowIVX0pkzV83GvpHe+GdH+r1uzqgn5YcmwMoEwGW
Oi5hhmlKnILXKNSyXCnUvUt9l6H7fPa7uZnvQCkusYmjcKNxT9mbRyaf5Bp5QM1EXYtBGohj6ImG
iZIZRK26jAK3vDdmEBELnOxHeSo6bYJf2eVQGvEi4E0vNa3oubDJTj6XJx7OtUVqX3gMo/qyHN2k
zuVCBu5N+/UXEEGAPOAA2NxnKZd0Jw/U6l4RjqVzR89CwZ13osIHOcDg3OTWvOs+YTFzMTu1Zm8r
PO9wKc/no2YJ2/hvVPNjsrrOt1omqD1wZdgzzQlwrr4ITXubFCK+u+qVfPFT7VDwhCb8ZiNB2VvU
T34d8HDQcjo3h/u/X8uFVtXSvtE3cyigL9ZK98MNwHIrb9JOb/urSOsKGnV70KGZ6OedJiFf4Uqm
991cOng8Dw+p5BoSpm9I1vj+GVP1xtEScWsNASZ3ErTH0cW20HbCDNe+bRpIo/1Bfzb8Q2fAmkkR
Ri9DY5bHgBLv02US4v+1eilC2FCejBdSmy932WJXDNA4nqyyrKf39dMzQ0EVIMNUdhCDLaYoEYO0
/6jLXceUHRVj4hLXxOeiVcTeZuQKOjLRQJALO1BcDXoXVxaNHlKIv2CaHdtvQ+sVvqyCBlxrw6y/
/vVVK/I0U6+142bIXu3VirJ8O5eltsazRH6hT5sjKMBusNF3dFyqFKOJ3Jv3JVWolM4HGIL6xkIX
Oj9icMiPzb1FIv3pA+HKe/WQcPeDkyOZFTSYtzJ37ArmjIWNHZAcAsVvsZNalUoFh7bgZgQUMZe1
3J8mQ5Qk3fQOwGivZiGQQvv7x39QO9kEJ12qL6dfUZbCQQ2MR/W2/Eo6WqbMeMMPD6KJdbnMMRaB
G1bj5KFOxXiJXpNWZv99TSQgbUFHFqyLW3bo50y/oSLHYNJ3iZ0qMOPgBoVFVwKbnTIpMp5glZtz
r2WZwLewhrXMwzlGClgB7Xh44MjyuUgIiaUsLWnz6nGrDoStu/uFtkHTjOFNkCvoLVulxqPIlWvL
UfiKpAeWiUiDR7Auc0TshFS5nreQsH6Gv9uvJ+ntt9oXwrRaWkKhDa+IA9m+c1La0IaokJqzpUwU
DYMQKyUwn5ugNz9kR+r2FOSslxZnffQhXU2MXWd7ZgJcKz5+II5LPKw8DcTMDCvMRpcBcgFdcT+4
BXRHY5lESQUKxBrK6Ib91HhJJsLL8t9lTxqdbIyBFOxAXzv4m8jPcHTkBWdz/Yt5yT8HnW9aNwwk
N091AVf3IqG+r1CTQwT4N6BfergauKuYCPxny/jqgOERKvNvEve97Ki3y+FAPwgkI4MsRnjrcVNw
+dWfzTpMonqGuKhEM1ITaOIKdRmHNvRqGn4yfZc9v/dZAKH78O5514YaAJFVwJHiujACN+2WaYDN
dHt7FHGgtSm2jdeNEplPbEheAZ1tOsW/E0ZiHGdNqnl3+mp40xhlJStLQjNiqYrNvU+RjoFbH3+S
LLmLokizLZvztVlGPu6IGmbUsLSy686kExJc1Dd+pck6kT+S3tQe3vCNKX5t12bAiWD7sRGGLzKt
NrPUvKZJV7WAITLHuw2eGumbR61W30HdefoSSJ1Rm87G2xfjdonbydjnGp45++6VM+QADYSLWq27
UDOI723athjl2AsTplZtrw8wsw4WI+0DzwN5Bulful7MNGVXdrajzeuhwSz/ovrzQ3QBBV8o2+Iy
39I3OV9tbcFrVDJ+m5MpW06rLJ/MOHOdZRdqEGq+syzj6yJPrBOPaahmdgz8UJVRLqFsHsF835d3
seG6JKiHQ5RAu4Xobu+8fLPt4+Sz4gHhbM2NKFfHe1rdTmwqEplMww7U2PetllgdWHGkHpC9UOLg
qOEnsGKPv5JcEmzXzwgvui3Y994uYci6zo51QGHmCsOLBNHCJQK+Ik/3xylpqTAlPezD6TC5fKx3
VkAdYTbVOos+x241TbawxtRbfxI0NfVr+gIgfUZoe5ENIJSsew/gLsHNzSKOQ7FipSa62aknCh3x
XQyc6qlWM1nGLAfFvJKqVEKXCFZox0aqNbATq9j6YHRjgTgxOiIIIDCvuc0PuiFok+Q29+gRL6sW
HtuZpxpkr5g0Gue8+nclUh6Wi7IQJMOCK0Mcom0HVzJIf/+jnz4Zsi3s41xBE3ew8/N9hV0pw1rp
Zxpjp+5oXsL7DVYw4tnuVtamXHPeCEvMsChptPQNHu6VX/N22hPVmx8Jy2A8MCjLFjiy3zRD4Lrz
FH5VlGvk3sJM/6hDTQWWNGPZxSocul9D4nwROauROOKtO0tP+HDz8xtFtVW/1WDcrs60+NJncfFc
7vzikBQ1IBBPXVSh7sSWtmpSbEQyzC6Itz/yoScpcsNuKWsL9bZdrV4n7I9Q5+vA4fN56ORDppXz
A6zsEoenmSYRcKxNMqV9YU7FzhPTll4D5FBAKnmFcSHSQKhdrqi70PZZbXHb4Lf8hX2Vcm2b1f5S
D5dSpKmwdNI7Bg+yeCCdX6w1kAk0/GYiFzF3TEAmNohW9i0L4mqPDOQh14jMxSVjF1H2n6OhT9Ex
WmWA7/5L1XzgNUtUat673i8fQfTDCJkEa0ss52Dc6BomdF7xk1/1ITO1cxF14gVnvA5G2M4cmvfI
q6c7FJXkadpU3lnSclZpQPXW6pm2RwG9pTtKIUXtriQSqH6sM15M/tB5XCQdllL6dViji7BfRZEp
NiTfBQ5uPsL0UYc85qlZDaYHXD7UHxHXCGyF0m0TySpo0DYGlW9lTcCTmhcaCCrqQbitHakxsoW+
mM82Atzi8BcelDJAx/HZFQcYTsFRJyHDSFHH/Mu43IlQQxqRv9kExwxSQmGaC6JyL1ycfBPco9B1
ZUwnFGd5y4RFXQI6uJlab1G4Jm4doiJZDrZaJ9Li0/A+Elz95t5mcFQMSCEzPk+mcfHifBLrqvYj
V4pcv1e6z0ZI4++4CgEgqHuVfpUxCvqo6dksNsNw7Gq/pcCBKE6h+fId3WXeU2klgpRzVJ98+zxJ
+uc1NGwcj60Dbyn1OXNPE9CMWzgHxOE7ihF9JCXJ5MvpI2BoPwG2ZV0uj1NLx6pQvnl8pntBXKgS
QfSel0ndrx7oJbDPFdk1oNR8NANPmLuaOzvII7gpRgkqAkm9/sw3/+y+Kk37cgA0ZUgkLE62n6tS
+30NN0tQopVFhpV+qWnf1873Ds3UInKcrzYKoMahpbnXDkS1v/h/hA8ppChJTv5zuY+BsvfnTFAi
Xv/ymAGPKtpvGLHnz0bU4+MPnmGgtun3PwI2d9U+ovQ76Qt+iLpr+eewClzcYjeqWNinjlGX41uI
G6nuHMlOO10TxFjgLmaB4KyJCufBjxJtyG8Tg/PTeWkPOFaXl4lA64WUzMkG7x5bU4LxvjKQi0Ka
HTBP0xbqIW13LnCVWbD9WuI8PhLWV/eVg2okvVX01o3fWGvGGoDtF9mgJI6ecGALrXJW13J7skOl
y8HrthO+PVx0fz8x+pMIaU/2FOY1qX3Pn72+ETz5ps5fcdJFsvtnLCBS7/5ZbYl3EHbX6mckpye3
Q2ZWdp1VHvThzJhqfeNyBSpUwLLGaXCzM9qsphupF2ccjilo5nOThez1kUuTqqzBqXbv38m6Ofvz
YJpo0HZnZpiyUbNlPWwahDJjvoOEfTyPMLsk2SbN5RrWnGl5RNJ3U1vjYQmpa743EHEA5l5cG68a
xmYZ/qvv4IJlVdvQ+aZ8oVBm26LBpvH3nmRhi9ydOOoRDqFppvyUxyj5XWwu6WHqOKmZDGT2Wspw
yNd1hL+XCAN6NjYF265FpTV3cEZ+XQluo2T+XLO77meVOLTV/3EvoVwFO7BcszPncTI07HZLtV1X
37VJTycfnwgIoJi8HC+q4fI44fY6tIl/VcRYEB+AhJPQgDRWvHF102AckZ38AcuMiQIPXQSmN/D7
YoU7S9xEjmROZb5l7cvM4nQm3x8/XC2sRTAQ9FQmleFc1HTNCnzMgE+HtggIpDiUjxA+/AZDJ2zG
0uuVmdwmJPpJYIfH7yBH6N9ywryUfaBQGU64ijj0+iNAtt1kQ5vcMb+me5T7/SZEb1WeZV2iNqRs
VRDZge/oX/KSWd9KENMEZo3nixjx4X/gPMckDXX1W92Ji7yp+/0/7XmXdOYQDTzpLPRDum48BQro
zEoidCFoK47QheDjK610zvpeEcbtbsBiBtkXgrhiPTaRnskf2tVyT/OwNSpB5Anq2tVWnf4Ar/2Z
BD3H5UjzZgt6c/sEPQVgLxc8DUwWmP9x/LS7fUrHiIm6jfU1cVr/N6DmmB+Doh9O0jDOMgZDj/CQ
mxdwIS0GsEVGytFiMCNU79A5GL/PcITAh4qdBJw9yv/hihZIsrXWlxIfVuvQm0FC3KztqiuEEcr7
XguQXlZGv5Pefa/Y11K/JYdF72lHHqxMCcqqHtYKqC/25DnjzBx6EG17buYr9f9eofditXG1BKpm
V2jUzht2nDdVcw/6e7IR/2MyysjWiMr7PJQA3uzJSkrX0n+Tx+jV1gaKydvrqFBci0REKV5VhSFB
cJoEybiqbJJT455QuLDk08k3QfoYL0F32kZPx8qImvnw+svMbldW5JZlY8cI9SbJE92S2rSfIheI
jzsptevPtrAE3xQZkZ3P6Aubbo4aUuUGJTp1HRTpO/ZIChETcBGHEmypGak8AZL+3C6r42aWDSLP
oeBGPSJA1ecEPfyxbRA8RyQnenm4yw5GPivC0UCcpD8YLAzZB/Lib/HDJH20LE1YzTXLVpLjrnLr
DYiOb2pkdv7OG0cw1sGBJ5sXix9fqJu7ZzsomdNyIP4Tbmkl5wI72qs4qh/YywLYgKEGVrfoEmjh
VXWqawO6oZOGP8fyBAF5tjkkRWdO1RBluyGy2Plcm/AvLncWckfpxWRb/QVayjtE8y6hUiKMzmHR
p+S3UjkPUoUfcyHDN+hum9hPhueTZys5sJE6rM9K74nsDn97xt+ic5YTB9RK19D/f4HozW4x2ITA
lsTm9ntY/Ucv0Vi6/92JGUJwmv1bv86my62pIJcgxufvmmkk512j6b5S5NsLh/70zDx/cgGum5Qg
fQKDlZzwxmWtk7xDSC7HLVMjtrC0LlcGR4jNGFK/FdK6+w3keUJgQgx+9iXLJs7btxB0g6u+J2Km
nCjYKG2nJZaxGk3ZmyPvVsCVJ0Wtmqn4aSvLt62Tm5dkSDg3KunPzeIIpKw6SuMRFlbEnsxt1W9s
6iDzIS7qE1DGQozQLF1o3846xMPOkBWhx1Cadcg/+WZDlxA+5z1CZ7OT7Z64SlHuFWzr2LcRdwcs
0I/JL0OYQ+zTEAZqapvuzRKE4GQb6Ikbf0+wcX3cpSEQq1oF5AcYTvrLkiwPxkMzsA4cYSzTz36W
UQykdZFgvi3zMSmF6lyvRSQ3dh5XFf4dPYhDjq7UAv0vrM7MeUvqYfqj1rBD9pHR0uuSg6WL1hp3
b+8tEwHI1a0MYWethlA74ISptSNDhYphSXr5OmwJWvyPwv7zRz/jMgADTXN2tTX174lCi6kGGP+Q
rtYHRp/0DIzqu2s2FU/MJnO12lTZY0xqwf4wfAuJnflBKVt8emz1ZE3t2wqO7svC7eFe7GETr8X2
/nYSN/V6auFd3Q69jvZ/OmwC6tmPHtye/xK3/xAdFbHC6aFrLLqW/Ze0m3GkQbNcabDbtael/8wj
tzcqc5+k8eTRuXSDeGiRpUoZfUkr2SklM5xqJ5IQyzevY57E+vyKPfP8tp2RTlUQYIwYY/w1nmv/
VCCjAqpZ+B+7Lm2VYfhqqA4+MDAztLXCM9g1GZKAA9tmJwtev5ORB8DPSBZwZkDwKnzaFyLE1RaO
Nu8jBmfJkHvjYBtnEtIfrgGd0PGjqf94jOh0NBvRvsj4DyVO//6+5KL8aD8mJmTtSjrFPl3u1pse
n4XTxFPCXwgLuV4Blv55h/IqmhSU3/aOOaveLAVlgqQysOkHWR3+gF8LTUMTP2yGmvzZNt0Ygu7P
4JBGzQRAh1/fJEbiM0Rczicz0x752owQWs1w3qRlLDwHurlI3yq5xUxk1RkB41s19yY32axz1kOb
Nmxb38t5HVex9GxnsgroD7zHQnHqLl2cjId+KtdQarhyHtcJze6UpeUtKarP60kD+O8wbxVHFvnZ
bYAWoK6YGZmgLwHzd4h9EYRcJy3TOUXD8DzNBD8jxRvBVZkmzEaSakIf9tZjFPorQYtQARzuikHx
1xwykDx9HMAkGWUBPVwwj5KJGTQoRgzILiu3xiFQUgSDfrJ1Kb5fae0CSCUzHjPABDzxclo4IL1Y
eW+pUtNCQmNhsrfNxDdcYeKMdP7xPUsRtM2MQVu/Bs3Ga/dUL0dSc+KIhAlCKrZdacaKZQEle2e8
TUu1YQkwyO3z/Gd8tu1Eo2DxG76cLpD4wxhlWsPdpT72QNvQP0RLHWZUXUNm+EG3/01pi+5PVEwo
kYTLK6zm9xXm9GkKGsTrEd/tA65YWr+swb/q6Fb+NvhMA1f8eQUPl5uD3nKK37SqhDEf9GyUAJVo
wvDFLxHO7wgkT5WuHMaq3ghtx6d5cz52hm/jrxwWmoglS/8u4zXKa8gLjvWphkau/JipBsqytJ0p
x+9nVUfJiUgG20VjTgwqv1BCn6Fy7CyNZ5fCakRqBXzMlTXuZ7C0lXQOC5oPEpEKMt7UfWnO0Qk1
VaZsX8iR/hBIF1wZLRlPzQyPmpZMTd0MKspq6R9V9B2uHKWY2o77snZottE2GeZYiS2CBZ8nyGSP
2FnWhTRlgiSlwvVy787Ymrh8yEgAUBweKMznftnrfresEWt0KQaOVCPGGiU6h8F3MpCGP4QLKPtg
OTXZFyZB29/7Pj2As+OaVxPQYuGO11B1h83lgTfXIEU9h3gAh0iMutBWuDcTUg7a/EvDYM7J4Y/k
BlovTyGiLANQlo5cw2GqmXlM3aPthZ58/IvzlRI65D6kJ5zpC7xlecNDfDEt9FgcIa0dpyIyiTM4
i/aJDHqRoiMIL7T/0roWo8/W0SRrNaSIMMSBnMOuU9xe+UlTz5MC7jEt253KdUsdGShufzmmtr3z
DF+/p5bZf2ol4mffR3u2MCOejMjcYO3uPoB/VvWc86wDlSP45A1t16GOV9Vt//5yK7fbm3p6SHET
YJ6Wa6C5PNv/XEPr1NeN92C59+BwsVJ43Czb2Pm0x9M3PmwEuECmiXXLk828+eWNVGCKi1AJdqKq
3S0qOCt1mPgOaRyJYBsVuNKC4jaH/fIwwJZzmMHQZlUj0A9KLUvNtxR8tDzzobZVlUoklT/6QuP/
3optISg0BViC5t/NnOlBkkm/U/XBdiw0DDs8zn/iGnZ2KYBhNODAFzlC7p05jcybZmrXXqIGApo4
zMllsd5d0tXsqXWnEw/XobDa6sOtgCaGjap6+TeRBkLpSas1yerS2AXHB102YOaejhbMYTwZ1iaZ
z5bn4r4GCoP7zHbPkiS3vagLDGFNXzp7ps1bAZvAQw0FNfb+iMgGDF7dSYHqKY8l8/b3D+0K3dJ4
MlxxhDbBIIoPkn5H6oS9MS+Zle/k36WkAFtmY85rrBqYLTrFSsyGjE2vTKXDjatx0E7fnmdD9y27
caR1CDXCV06dtlhBSdTyr6UmgrG4evVzhwPlxB/7il1+HQR0fSApJzMcqdvu6NmYfQUL55Kw8h8P
LJ535cXkBS0poq+U3FLgJiU71WEWRVAipl+6os3Du56tSfbbWYy28iau0g7FGLdjPoFgPXqSDAj6
uXDpwQ0GniWeUQxfvThtM118u4qIqE/w2PL34WrKmEoCzAdvsrhFj0qQ0W14W7DAffFz6esUJZvd
ATxTcJ2XBNsGmMg4vQE5lmEE6jcobaVO7phLH7gx13ng5nN4FSBcDPXi5Nfj7FhVbbvnMupEWTdg
CSzMZkpeovYbrL42nb7ARCGq0BCmIhNGYcY8r8UDvfHUrKm6W+HB2AoYdH/e7euNhCTuzv5bExSL
Cm/6ZnZ4UbKAmTuN79OUTyAEt0bCcHGdhpWfeiipejymUw5xgZNZyCTGFsQZOZikzS/uVKjxpXrS
PybhiZ2fnT2NGj2IYsjompQqgYCqbwUBeq/BWsPht7aEt8Nq6LxV54nUmIZKSLCvbfzVHxUi2SyB
/NmLFR8mDXVmnoguXtzi/HGVDI3UqpS17jBpmJbB6HFC+UxyXI86OH+fgdl/SHlNQ4OiPKKCbbZR
/kktAfnErBWCk2pYxyvnmH/XAX7XJ8VRU7CeK18yrPNvwmuXAk095DKeHe7/9CvV8oGEiQep6/Cg
iDSdK9CXcRAwn/M2JmIYv1dQ8pkz83pk4DHUg2I2As3Qaw8azT6by4qNV5zGvB/oCN10Ks/7Cnxc
/AbzVRCWGz6JUKRf8y58IzpdgxUbsmmVSaDJmwtW1XhxCiEEfdzdU/LGbdRKrTPfSQoBdq3j+1Q2
/wFnrRf5nTbBOIcuy/IZbITssnr+puksvBJHsiC/D5IoUurFWPPlBSudtHQSsrb3/ttWPZn7WY+G
TJVXRQKstUtQqd0EcCCPNU+I8raPeCJQkyCXiI0cGjzH7XLXHGzOrLVKIjuw9XbeNH3oOoU4kn0O
gN/x6iNdjsjvnT4CgNzEHO5yGq4wYdNqudhRh7Y1sF76ip/tSbINAyEO4Et73nDi03tMIFvoISsM
jv57vQkflld89ZAB0BJOH5BJljtX6nL8rDQ8yDQlNXLNdZBMCtzliI+1O79kRPPY4S0clAY7BNZx
JLFSY7BP1AZB0WI1pmtV6MhvlWp7wp5v4PndU2xIZaeEO4M2Luw/hHx0tSR9FzZoaFs/pxJBUC5D
H5adlElx5PaWjl+o07wGs+0DxCDTNBeB3I9uBoKjc4wINrUJC0hk3+CLlWzbrq51GKkEkBdgb1OC
Nuu+NvErxHnmF1S6HQyPq8rK5o607X+NUBW4DxN8F4HuZwOs/171k47LCCKMVbkzL5qwW3QUQPm1
c9OIdhb/eRdoqn5VytwVUHMHxA8WzT7u3rHJZu/tnCwVnjiIQTLEth04ad6KaMaX6Z1ek36jbpUE
jPI5dUC/VK2Us9gxKN6dVzBt04iyE2KAqX3Vwkid5cTFRRu+bky6L8NY3Ussj0acx7MhxghpaP37
sGhN1Je4vxX5pPKds5UCkYD5TGfS7AIQ9Gm8aFJUYEM78IzdPFoCMl1ZLeIFhFa/QeRE/hw0HH7/
tcJ25rzx6fhzBFBmLorvd7yyvCcqHC6KzlO8FBLtv5J8a2kKTmo6Vho/jUfMHUl0EKbiqULL7uYT
rk6dC3UfwEb8G/D6FD8sLf+BtXaLncQzhZVviOOEz5QfYIYEiRL0OiarUVpxs9kHNtid0zj231OW
bcqfbiMcmqynlDH15frQz2rrl+JQ+96HAcPpN9cL1OTv1YAtCGfs6985ALLU7O9L2WZVuzshbRyr
zceCz6JQJ3JRFJZBuB6O83Yx3BNEj7SYzVmdyrxAjYFOVf0f7TVPnWoSZO4KD01fSnuYFanv6CuY
R5QWmmt74M9qYeHk3mGCL72DfteL1/hGB976x3NOdXb9o/5aOI6e1VfY4Ji2TnehxYBICCl8ROGN
puqX7WD2hozgIo2LpI7p9YCNQSK+S53ouc0cnUCYQHx28ryauH6PXoI8C8c7p7OVpBJlk0F+WPFe
/rSHeGLz+6LXDtq1Ozf0Ajs1RUY4tcTjDQbqF9TMEM4SLwzBn9tf/r/vBOfc9NN+Dw1FT7WGsMBi
Dkiyhy7guWOAGLTWJQSPaeXoHJ7YR0f4bOqbHZ+ZtmmNRoAd20Y13M+WvXwj3y5/4Pk24yxe6oc/
A1YdOvBNKFiouMfBbp0mmiIQmN3Bt1E4MvUstPC/btQoQu63Dpgwh0D2uk6yKunPNuHKsj4YMtUd
8nun2X5dYqc9luGwz2laLjyuuHv9ZNEeNSbG3VvKCBi6EpSGW5xSIrztbOmTtyzg78WHZRbLbayn
3Zi5qID8QDaQyiMkCGKx1JYl5I7oEDQXzeZrT8MFncZCZjDLi5fjJwLzm72rTG5Eol5Iz5I1tOBj
1BX/EkeDk9jsoklSp/EtN5tPc1eOMzJq6qSTgl9Hbie12/j+Lsd0K20grbkvPGLcqcP5gu6WTEnR
0Xj8o4fjsTGxrerIKW5gw4d1kGcy+TwmFKlLNbh6pLNNUdlNP9aUJcAEgC76ivDf2OR86RmMFj4y
aAp27JWwzElwcZ6oRe+Y1UVQhM3FZEomC7IRV1fjxm+vBU7SzXu2OnCsaJ1hGXnOAm9xDODXe2UT
PaJF+i0e53L0FRiKWT59OU4GSvqJzkXi2AkOk5eKiXgonwlgA4cLq2XfPNidfxZjO6jKMcPHzsrY
6PkuycUv5qqr49F3nE+zrW7/P2FTRg2NOkG4DbO1iJjEKhSEQgvk3hLu5DfaT4l2NRIQ/Gy/gnAD
UPGT9SlE1GZ1c0kBENBg4VjAp9J6i43pdlYiGUHH1IRAeO0DILEmpGJnzGLblyn2jaCF5i8r+8ur
8ezDsuHnsAXe+bL49culGDjoCX7gtFFJN+v2KlD5QKsQ9DTBVQv78GTy9p743W9Y4WiWLJ0sS7jY
RKPm0YwxeRbFhh0mfmvd0TPUTrJdgWHP3sLqVKWLWjZmtiwXXF0eFi5TlQy0OyOtQP7YA3SHIuRp
AkZmeCzthZiRttJ0l1k1QCmjZCzNYMH+JLhXpj769aOywPHBzPWaKTWV9sitJyhfztvQLjOAnn24
DoJtrZNB338ZeuuMuVP43G1g3MjAOiQid9ItWScCyXK2P0tgA4bcK7IjE998ypmX7XgE7CFo70Qa
NNHaPA1oreQ6HW2FfqKcJhufGDI+/6ZBrTxrYJ2f62ODQAjK0Xshw0mZuS87TA2pRmj6odLIWRz7
mlnW8o8nK5NK9mOJnoCumGrDOws/Pu02lwWIYt2aAwSo1ILI297/3+ulqzxUeZ/kJu09vIfR4WI2
lBGcQ9qNDtl6XVgWxxRRjEsI6LAF3NsuQQsFT1X9s1rd+qVHVVrujXl+cB0SR3p+3Bo/1cpa5k6V
jIRXvHonRcCh7iFhKwvsTrewRGtFRzSgEI3o15vxtCeCosTwKAXW8ZHixNSdO2m7XVQemZoB08Mj
xYNK6fcrrPusl9JYcCvRm8f/v2owkgFVigEQkRgVPi8xoJPmwEr8vSgKTDVUEcSQTCkvC6x898q+
aks6FcdH2GfZ2tp3nC+3yCM8bIUIcn538A2F7M2sqZfWpI9mj3H/Kbx8v3csM2UrdRRwfToaJc7T
Ry/+e1vIaBfi4SuLWYoEQm0D0bP9OzFkPnaTzjCcrj7vnk2jPDcR69TRr4d6BUSEfC5Drh5nb6+v
dvij2wW26R+rX7pbh3U3j5FSo6i/SGj8umuZqvRWIrK8kaX/ocw27fJ6d+9tMONI10FGP3Nx5zT9
NBI7jLkucvNJ217IAvd5J2wRKnb4NXjcnXH6MpSzYWuMBN852ZkZkgcdxQ9sfN8FM4owDE+WBykg
P8KHJ4SkCnOhOh+mVuG1xBRJQyZsJHaDrelH12ueMGr8tt0LsTgu9j5VwHd2gozAYva2wbxvbL2G
V4TtdkyQSUPRWiIEFzYEh487L9E/vcnaAIVdr5F2vLfCGlKXHjrkiYu6AffMTJeI49d/RdwdzOGq
r6ZJEIvWT3DFxcpDQTN0ZV7aRJ2xjSzTXMrz6uaReNicbb1DBgPNR2D+L6hW5qBmGaJjb/WWCeyD
iCrV8Rcg24squHCVvTqjv/le7EU3+yX+hpBInl4BtqkBHGHnAY+UkxvyUykYb0jkEm/5M9comTJd
VriHXO9GdECy5LZTerQgoRedvawWybW3tmsAJOub4i0KwI8NHYJYAM0UTQDg1vu7HMRUi+Wa2JPB
GiSzHWHbTdRqDc+vn6wzM4/zV03ccHIMbfUjRbydzjYfJReaAlXMqRhZIjht7NEPTnJc2vSkGYTJ
xRtmUUWb2p0xLoDz7oe2xs4TpLs7GEm01mTG8JA05WyDjad7sJ8dTR2IrO/WzsLjEJwSE2xANMjx
TJm/whuo0sfvlpy93Mx2PUm0Ta8usGvP7bbtYSS9ZPhz1grLIS5iLbP7lTJ0+25QU//bl9YUNCV7
ebfkGNVVtRZjw/wedWbo49FM/Fon6+HPCuach2fn/u5hL1mkkUoW4O9J4DnCnCDf6OpXMgA6LB2H
sPfDu2VFBoaOk1VeBokYG8Ag5CDcTEEJMQBFByOGgOT7a94mtOyiWT20FZEGtLGwzASYHlEeotzL
Q8gWgFw3vW47onu6drtGqGkA8TYlU+WjitMxWceVkM1Q+fftI4Fs5oAIVGJj1zPqzl3YH3I6Ytl6
tKWIPC9BSHIiogOIlRfbeO/l27aKY5cmB20/LWbMoT8AQpJTgKZeLvWGdCiKgm5BPSXtIFScOmku
+9Xhl9HAa9PADuaN5XQZ2sZU5UROBVvn6l8VjP/h67qawwkEUbONVylN84B/Gy9LMTK3TrOGLADv
FO2m5OmCv8Fr2yDbvVLEbwRumeM4bX+8qVqo5SHU4lx6zKieXMucTCvSPJGEDRNANMRreUJoZSVV
Yqjp0MkwGFd7uHbkiAl9PBW3EAOBVVcAYq29EYJ8trputMXoFnQMIZ0CRLZX53ljcMJOFqudwAvO
IkJ4xwlI3Zb3dL2KehvKRMNJMECMqubq/3J6vAM1/0vRpFGhd+GagdrMwW0Ura4dB82WNkjVmXnQ
cZ6sNDa2yx67WYmoClp3A7XCO62oU7Bmu6q5aA4g9x4yizmFBjzvS0seWy9g/wK5Ag+W6hlFlOEv
f3j9+tdAgfli+/gSaS/WHGYnke6UnCmjfqfLHqx3xsO1HiShGRkrhV4r/KLw0obX0+nOUPOENvEF
yu5Bp3LJNtv8eJy5ijL2L7HpJqt37Otj1MxrY54Uj77S3BUVksqzct2Yujh1Rq7CVzsFp8jUfpRi
rqT7I1It4imUE8IHDhgRsSyLXYT3kyEofzsLp/Xvg4rJQ80Xb3KZR3fl+uPHN9BI2QJOh1qM2DEe
GRrYg03jSEFrrepqkxC2cOxLC9r4hZt+7WNCIbEltBQs60YDivMUSYjA3izBe3zeUey94lDOXbpW
lI0FgxSm1f/2UCAhAAs+50MgTwsjkYcI3QgP78nuQg7equ1tIBVJXLEsVeGT48PSGubpwU/gAXGq
dSR1ou2NwtAy3QWoFLxEF7+amU5ns9BZFAxap51p2dRO9RFHgQNPIdKA7DrC7Epphv2FY+4jRTNA
/ojGpxxPD0F7Y/NXPRRECyh4DcLugqdYWVPNyC3EqBtMiaAk7xVM59AypgieIPCooxg79XPTfci9
6YxibBuN0iuSSQWYPZcwPpremuFOpO/716Eju4vZ4ZqVL7Mlb+jxDAtB5mw1JLuIEN5yANdcoBxJ
zjKJEuHf1w2fejascLQXbJWoEWHSpAPNx6oDCGmyOiZcHZsYGKwtBp7dQ1YEdd7/tb93NWzCQIj4
oUvs85WcLmQ8ThB85HaIU0BaMlwco35XUqRAjmn6Yxe1RsblnvtaPCapQEVlkx/UvgQXVqGksCQJ
Pp3AecyH2DFdixe/R6fZN8dx8MNKdElUSC2lB99RfkK1D2S/DvcUyJawu4vm+SyDL2w3oBKfHBPw
R78aa4memum0OXKdLTne5/iW5LXMFMZGurUfZzJug9viyx/ZWrsKXgl40M1u5Iord5+36ERODP/g
9P+K//I6eLMPZvZQJ0RbiN83seyOVEUWT0wYidTCrF83Q5KDnNUQ/h1rT5fupf6Quj+iKRNm+Q48
BqO/LvpMu6NkDZkVCM8y44b+vdt+KNe0M7uHbacaCQXi+xLDVatNNwq+FAk0Eu38IHnXEHAA+jT7
5UPy+5attjxYSxrzn/pQjgfKeHr2yxlxqw3I1fp0H8W0+L4ZIXR9KHKMj02NQqB0lgRpGN5e46uW
pETFs/fu6NFlJbTEkXJxcPZM80mh7IeaALcFCBRPny3sw3eHidQAtWWP/XkILSf3CH8TiW3WICo7
eXVuvKXQmUVpg1a+AgDkLEHw9FNwH7z/mhWaJ8v0uO2gIFt3WieXYamCKJqVqu9a2lbrwa11pI8e
5AJLL4d1KdhiERz22/0Iy8yFXok3TPn7wS+nSYARNwx1h/V2zXM5fr+lsGq1QoKSw9APo2zGoBFz
H+64qZhPVneERGZ3Xe4Eww5ojtJNz34Aweu7YpKk9xshN/vCBOxZuy5NDkmw+r1ZT09sf/ymf/Uc
rcBPsXvs35ymtEJzacdAiQGJMXkVkYpxvZZkNhrXSOExh16V0NXZa7istU41TCjMfDmlyPbpgpWS
E0mzF1Dzs/egZG5bub6wbuZUyUQEUj2GzjFJbOuAvbtkkJdUkPPJUoPOx6wOFcxieq1z0ROp/vwZ
diPpEn7HiKBjsA108Rfnsh3A0BjDkSEWBYB4fHbRawxO5fQWAQFym+daY2RiZCh7F5ZQjaH5J4cO
7PYvd7BQNFZ1lrFbS8LkAhkxdKvqZ/ZA23l5F8iZndf1wRvDyvaWDBP4dLmQ6cuNKljDir5OTHnX
570CMhSHbd5e546PPuvrZg9mgT38cHoX310qcH53riAfVG99LB8PjTvCrjAJTkBBLFqk0i6JVV0D
Lwz3jromz2TfxhU13OWHvY6o/Qk5YnuNjUVFWSwMO0lJtiNbfRqF8fVByBwVCY8p2+g4FHmk035g
2/Vzs346i/o4tjbVAp55du93TXMULIbsPsfiTzoAqE+JWfMiephzSQIlEKKBRTciBSbSA2YWdW8u
ZK/M/0LPLb91o+6nY36fqzPUiRKPmi1ppyRGgWld8tMKUSCQ3qp7JL77carfd0xFzWG87zoV9T4Z
tLbI/m3bXdDpmgg1RvkYMONodSuR92uC4H3obJNTIVCAx2//KxiFEqoJ6UH0XSmY1c3HuGjSfu8J
rxnaY5Sup5Yl9qZZSY6mRMkPtEjiDkU/+h6PR3y/Mt8XIrJaM4P7eSDhrXcFG/1yuEWzvJ+tyjT7
9cIeR6DIcJZU6n3HZT/616m0QF2hDU26lL7j+DMkyw4sJOksJMdJ5CkHKRgQSEzte7XflNWcgFfF
0QnLCEgyxcsVTfy3u61DLj8oYN0dH01zlohqheyAKSjdtw/lHQe2So711eo1CWZTNz70QM0xuc61
HxAxrR96lFnduBp56mw0IGc/rI30vAPlGBB2x6neazvU9lengv2PWEwnoOhTjfAecmbgwQbptHk9
hpMOoHmQ0b72Tg4j+QTDZNMk8erh3QGSQfgaDd89QOzoPOOPBZ0snGrABcHTy+ZZ6nkY+RfYa6R9
MwdNIEfHXkrMsHCNO8wONt0cYp2THz5MsgePdtn5iHYArqysIV1uY+dvXimG3rkGDHR+UvFjBvYU
z2TB29RsU+cT5WMnZb+CRSypiafio2YC0hV92zDkn+3i94Otc3gCU+Qd+tqpdxMElYO2Y0guUi50
0wJjfUgvWmj+9F3OoedepEGy9SsNYIIOkkDoAAPOy9o76lZBT+OQobvU/IeLa7OoadKQB8w5bMIG
VnqfAb/IRFnC0npVsOuDCXUNGXGkKLyWpCugHeyw6m0nPMb0lNS4n6f+u2fH4oKdkrTUoiDxRRat
Eev2rUGICVXK7CDOcPAnhSfVPYwEfJ1HgPioeBBfT6AtKZTHq7rmNQKvC+ZfZXPo5QjKAPzM2pb+
kfzQKkGkWcrSR9O5l9tlmo54TIeos6uJIKEcwD82vGUKegQt0bews0eIxq2D6udGAsez/Q+uL00V
8BZJOkXoOfUjvzMPVBGwgl+NumrhLfsX/tdUc6/+R5/WybKp3CK1YgAss190v5oQemV58NfLZLqX
uIrgci1fVs5RtEnGFUS19MPeqs6XTdIn85uEbABoXEq+jYGkijAG1cgFcog86Eii6XVH9Z6ZgZXG
GGI2lQJ5mYQUxdS++B00MXIl0l3ce6kjgkjGpOIy3PrnCEhud9Huw6olcwfi9rulPSD4PMvUBq/f
Y4govK7qgylX4pXItaMVXOb37VQ4QLjiV4dqZ+qzKuHw7VnJH5zJZuCd2bog8mZmByY1mHHttu9D
Dd1gpxLgJovy+dJQcpFII/nueXbr1g6PvZlW0Gm3Lgrdu4zpHDoRB8dgolL5gt9fkry3b8iqBOOm
BUMfLdRhViWacZ0ce+79E5mfduDz9PyJJAih+eTvjTgnrN4VNe2X1Bd0ZnfleoQ82MaqH+tMPLp7
y7p5s/0nkHPEeryYOfjG2VYg9n1DocYsNKemd3mIAM89Sy2Zf5QMPw2RCmLk6eNcImLXoWlk899L
vAi8gnycG4p+4wJ9/SoUJUqrgFM/9WUo1ZaBjy5qMB8sRN6x2R9e15LpKiRG5hU4ZKW85Ii8xZIv
+Ow8yVinZJhDiCBpwcJyLmpx93D7mUQS9K5Fwsoe+ureSaFklYM0+SoyA+akW35xaTTqVuWQLZu8
F7bb7X/X1Leb0WV6EMjxtHU4C28Y/A13DnET6JEc1Qj8/pMoAL5wbBfDev3V2yE9GPA1FR9Mjv8m
AzEwRL29VxaPg7hiSrmR63TqTqQMVYVn89Yb2JlV4QbzVnORdogUWclBuqd0h2zWRrAlHML1kbjJ
gmC0x7jU0vGA/GOWwL7Hi3UtYxd5p4d4WpUNpCM0GAyk9hZWLge5EKboW9orN7cSzFD5jSGxrdwy
k9PIsXbnHtf6UAUt3yzNcqQMsBZvz4JArNJRikhEiaXATfR9WBTEhQmu8oI4YHBzicHtNzJYn73Y
A8I76CgUaesH5glxgbLX5Q96l2PUEbLcUnhraOJKrt9yenG98BnrTPRfoYlax4c2knazxjuwgB8f
oOfU3FyWI3YKZ0t4HlCW5k9cJp0xI3WkDsh3Zf+iXVt4PPh9BmgjYWcGDNe4QSbWRhj35o6s7hF/
Y8nh7JY1wy7oCRC54tdgTUfLxghFHOvF+PCPuXD07q2p/QalEuJVA2334CwofFvFoQ85EW5/0TVB
RZ8Aeik4MbRCdpOoVqIziiV2YTivZHfO9HRcVF34ytBjdoMbogc0t4UgIM3Y7OcPLj3aTyDnCQf1
sBcPY8dJaPup7+QtRu4xTzaOLA347Nz0sTBkJHU9ABaCrmBw609vTRlCsf30j+SYquUiOCQvgh2o
r7VsOmPf1hdMN8smqWBayoAUJxH3c8tEG6Yh/VcCS5wHXbR6IxQKaVfjh7g4r1Qi0GxhPXpYMGuG
zXQ2x6VkrElpc6bkxA6CG9nGbu0GUkVQAG4vg98ZTYumhoM7ccSXN3L3MtHU4Q3M8B17qsCbtePN
VAD43xI7REVGXAsmOlXVMID7oOWuSm1C4TFixeUh99rUkkgX9rJX+g9Cgvz6CHycZ5H2nVstHT7z
IPSFOaFpMXQNxf2br+BKOm55p3FArlKEcQ7XWyvP8XlS0XEM9QuqswcmwgNaGCnS8TYTfO8YtwrU
Tgstxxs4UbkJq/1T1sRAEY2VidUu1pwx2QNAVBVAr6SC+vMLsM+rfKHW1ed/COFfjsI24IEBSQHD
ghPpDwFDD2cHDV8O/Gf5PBsjmKAekT5hmwAp9pn+n0GnDINUGgz1bQLzn9lGXyZljJK013nk02fs
9eMvV/uVlbK3Jqm9U3TBJqkjt+DH5lcqC2mff/V6ushOCFQDInesFG15U+hdTFCx9VBQX/b/EWKm
z2Eam7Nq1d4CxgMfP0zF4KCMPP6DrovMXiPrsGPC6b9zFmRDACSZfMu+oCWYrnnIbj1AUEC+vPBC
9gHn6PEVQE2PtnuFaRiBnjjC/PjctZ1AaMURYGhZ4Srqn8gkFX7zZc8Prj+SalMEiYVGk4sfTMh2
tknY/NpPERO3YU4iuaIpUdmcqd1nvIzHOW6T8NT3vwvJKptKnaeCS13L5vmYHEkAmaF1fIRLTANc
tPQcBY+KbG5Mimi9lvXc+QbejjirjPOxh6eeLAor1q/2wlJ6o0QkuL+8tiMHFWf1sjfDoJtTn48T
Xleb9TryQPHl+A4zWzdVmBX4EaxyEKQLgnppovS3tDCk2FVBnlo4Ti9n8IHMEZ0S0VvX6/w5JfwO
INWOMLsKtJ8N9X9ixBgsvh3j75JImlsXOZcQRfYqcImMFHl+MQaR1fDaAwAIkjfQvgOykAMHNotN
21ddFc18yWkmtGuQoY9P9CsUONJYFOkP383XCDe8dabvhP2WgnsE2Z8F8DtUA9yh+8zJPQEytTHI
N0p/YMO8SYcoYcZla4qRgqam9cPicBTXStbFWWebxWbdlF+wQKI5dwa/TOatBGOQpy5M5b986k9I
bHNGmpSCNYawX7HWNCklE3M4Nig8r22BPtlcF/RJalgdMElfg/VSuyXbaq0AV2gergTxB/xhdxW0
Er5p5gaK2AQ3Ci4tIoAOdMh5oqqYBOYVOqy24HxCTwaYfvt5tZhWr44vVWNeTF/bLxM6vEeK15GG
/aAGqm0nQU6ixT8z9FHc3xKu/4ohtYRfLHyJ37JzGcUoaTpcv3QOHQal23wW0xNIRVQxk25veeSQ
8B2xE/+wikVmb89UU3uytUUccv4u9paYOTGgoYb791qubOBc1xlvx0GamYW+tV4cmPROUiF0tmtt
6+MZDi7QA4Cgt2Uxuw2/N2fQTL7LN/MJj2fkaOdpPbzSGhegdALA6OsPgLF2/FoXCjeoZ6FUVP+Z
qzV3LM+kJx8JS6VZ/PN/2nNKY5dVY1mlG5cSrscJl7esZ8su5kP1ZFKIFGyil2wis8EnGxSMOeD3
VCE1ekb3nrClAKn3wkNcc6iw45yzxqw7truQN6CsjpLGRnIcpOt/+1dnEV7H1Gegj7Hy7P5Mi6eG
PPphqM8Ta0C/IXN73OrbR3G5K5Jaxnw+Oa4iXoaTBQrwKXaKFZSLvaaqIfB6payqHMubCwyVfrym
BvheWBQQgCgOJBWSioH5fhAz6yRXZPMk8TIRjDHTRcVguanyqYQ3u5weSLyZCiy03P1DMFdEu8uK
WpaGda8n9wKcio5wlRpDYlQC4z4lndHIMquXyrdjrtZCV3/Ugl1CZmACwgIf4z3dO9RCyM6y09+D
SwuPxCxpFApASqSc3wXMVTpqtLq9BHyCnIqFQqeNu+Ai7Y5GLE9u4HP3SrRf3GlqX8QxONdZDqBP
L2qPOzlqvOYKPucuNeTkUS2gA94jjkIROcSBffrcXctTcwFbiH7Ii7Iafga8BQjZtfig0UEeNDRv
TIjIJR4QcZE8kSJYlFPwIh6zur5P/C7QQFRewKP4jLJWzPiLLANPYlErzSGjR4rGn7J0OxaR6RMB
17p6C9O1BIXpYBR5YPRNC5U10sGkCs7EQat/44GNedYfwCS3aL4iZWzCol4LuEEItxKulKsbGnn6
q3HTA2fmh+QfJ+NXIZmJP+OKv2PKwVnuURSdzlnJ9YLiir95TgFJc7zo1Cue1ib8DIeUCvQ/JKpd
fFAeYRlqlWTjrtKhLe9tEQEoze0G33scBuTTTy6qdcQyaujIITUKQztT9OIeDJm9EJKZFTbLJlgb
5s5Vz5xrpFPYnM/WMytns3cwt75LXgP1IAtJVrOW5Wrmx+nriZ1H38+Cwo7zJbdqyNHZaId03n7a
GDu0wrdOVrZw+QHEEy5nOxvnW2RCZjHOJQIXHsMQXYM8FU1dzpBN+nYNfx0nKi3sF57KtiVQpMZN
QbunehckJxn+KTL4ZxY9U4N9yhfFYgk6R2kieWOdO1Gn8KD3pgV66/yIYK6eN+C5jQ+DT2GeRlDS
e3cz98ocLpvTiAMH/h3PtusZlhZ/e+VUn7JIu/e7OPC8sDYFX7LI6uwDr6gt3wQddCPoo+ae7x0o
ObpwgGZVb19UBcEIgNsKMNE6fNgx21QK/UEPgzm/rhqDqwKPIncVfRPFr2TVszw8esZwU4MpQvD2
zvQGRulTrIPZj6RU6vZGn8hMrIDm/4ChIhXoqFDoOL4wWodbTOUwR8fpg24v8MH7N64GJ2P/rr+H
56/USjSIONG3bdAO1+1OzO3XLxgHttjG+mFxj+yTX5vCeZ0s/Y8d3R1VLNT9pCsk8KxzvpgBz9rA
PrXbwIM3yPbu1rM55bOPFI63WFSjKi8YnfpIc9o5SQscZurG+H6PJTdKQv/SwtNbvT/ncr5nUTOm
Qe2jKCF6jK2c0hoNYYUaU/YNNeyGUb4KIyZOwM2SFeQtEkKDAlUufWbKCj1CLBxgfRX3QS+kF91d
K88VaoK0lhrFCa/NWEhwSPjzNT6OaZQ0kXDMecEnnk2jyN9NnLLhlvKJBmAiSJ/t4GrjBJsCQANk
ifqSmZbLLJ0hIhP7MLy1m1Gb/y95SxNeQGsuo/7o2IYx/R7vv2lFxr+q9GvmPW40qmnBP9bzxP7f
e1peeFVuQhYG/kdX2tH7Tf55O4yZlLkrbCf+brIqB9EURxE9yFel+UusDMDyasdO0SVKqqsl4Sqk
vuBbIVi8LkbTGavzAsmdely7o/Ier9w30Wo3evKa6Y8iY5Fll8tbezcV7LXlCyVyP+msKOLmqvRQ
TBN3Y5B1NRrJLmsYNJgslfZ60wQdp2RFdOLeC3pjel/Y+2CqRbFEfX677ehbOC1lS0Oo1MEngJTz
8joBCNKnw6+5TVowPNnQ/Ey2NE4UhZODsYTd8aUFWX5j+K9zaETkhjE8CHGUKwBLyU/LW3nvmlo4
K/CD6cOAdu9v1VQPxVkaNh8jhEIzfsWL/qFHfHDWd/l99JNS+Qr/QrSPRxj+Lw68nfVLj7tzOlL5
b39E4DParDXG7MrtdPgE9OMD5kmZWax3sK7H62II+i3Ev4nzHxijRRqDemkpBE2OG3jvGctLbssr
6SnGz9rt4/4iXru9FeUvGUMYEVKIKex785+iCFhxMeO6KR4v453ezvcA3oEe0bqf4nQEimq8Upgt
hbD+g8UM4LTGVinzQS1wWenK21SnVZ2QxUlcZBOaDo6XfUpxmjYmgd6QNjChVKFpbwDEMFZOtA/e
AWvzrK7Rhc8aOz/n0zEcsjfo20/vRcocSrQ2ROGAc3zztPaKjwpNtNi9UeerUwCejId5Gr1EMTfo
j+T4MhnZiQOWPSlWmQXcGxYLdHnNQaToKEW83IEBvaaDdD7I7scsxa+0+CjGpKwuKFuerCj2xKtL
hettEXHedbhyz/6k2/gZDn0BvIUi+mupf21p+RB8agf7ojFGcLX4rGXXHQpMuP1MWiIh8Q4ry1Jk
+0CJGZSmRgllMZCzFpcmz2X8vHGHxkN0/ZjK4pSYVTAizT7AevqaQr4htEgm4dIfhov7OvBN6gzS
D8v9DoZX42i9yaVDszNwoGFH0m3L62/uels6x5mBr5q4J5srrEX3W2h/1IiS64JSVRiO2oYxUeCj
A0fUuGl4rr/3NbmSbJLEsv23qUlKkXqGWJqn/c1ICG4AznkW668c8Am0iraQCXMSNS4PE+qqr5pU
AvcQmtG9ES8MKnN5Vy8TrQLCWB9VyPzv99eCkMtCyxh71xWienhAThtcgts0SUguzcFts72iFhH3
f+bjo9kZOHMneuIgGCsAkQDwuKzioDrTBP7ZVlUcINw7Y4GS+d8t2LAEu1JZE5wxg/S5EhtCFVc2
AYUI9IregYJW0TkC5Z8hTRYKK2AlFsccxp7aEJrJJ5jDzTvMuQvVkMrCnLj8y7VEE2vd5V6srmmL
oXlnZYEV2aATSosXZlnYvFrO/ycmg1E+x2UMJwhMnm8+coYblu8IPyFo1YtI0YISFTTaHDrq6pat
3ugdVY6kn4AAe99hjAsor2zQfLwCzoGqYw8Ny1MbjP9XfFwTUP/whMeuWjuHw4LDwnMoaXlz+hhg
hqgFLOWhPJVnMYL/+E1uuZSA4zr1cy/YXnq/2iWMlU6nxe8+xIXv/CFg4oJTS0v5EgCTc7/ZRfLN
fRk1BnxF6lBFkRHyxeORar9c34775S9GChExzln22Y1d5dmtwA6xXfFdj2FqyIDFSi3SpK7jFF0A
4fL0SA0AXF88mo+H69Am1HiczBdU5xxATEErbld55AxH+hSbQV6bo06lKGYODFD/ANjnQYAXLy5Y
16Pj78k3uIl04MW/rEqJuLasp+x2nxojUAYTgoilfQbMhziz8c3zYBbO2BdwI7ZSoDvGCXwzNHdn
6YmA7wBg7+MZZKI9pX20+l1WLa7iK3TXkjK9FMRROkN1FbH3otIRpqmbMrBajEQthYPK8coO8CfD
WC+Qmo10H9kcK8MrOIllQ1+5M0s6IzvCBfTagdYx4wo2Y2Nc1zOhzEixMUtgfxFnI3IXewTg/f6j
A3lNGLMV7JNkbsU0cKpfkfJpsd2RCKyWxvCHPx6g9LH+TgYaOl6VLbCI/kEBt5IaSQgTP9osrarD
Xx6cCvt6Cfh4dd6+lPlVtMZyEWVehXIKlOBRI3mH40FXP7ouJkdnAy7M+/Eti2+QIfDb5k/fQknp
CTOzl8XyRtyqGeZEcrNYLJPQe7IzobE4co5OL2XxVYgpWl5USfCDAosH7xql3BAIcx5bxBEqx37e
WFCSTuYY1l8m21oPf8/8ORe0Z3wAV24+3o+Klrk6Yvpyd2nDw0/9OOOTROyykzKxnFHhNLBwt31c
rIGQUCnoCi5U5K4hWvZe237fHt8PLJ+mb4BY11Q+6ys+aktDPO5XgFlIQlSfdMaVQcZSMQKcbAnq
PxsPaydtyizC69xFRA9Dde9dYChIEolihxLa7LrGpKm+e6akCIJ3Urb3YK+vuDUFnKN5AeVnJxLD
XmHYjGybzpKSzriyAahTofU4P0y6cmjSiHox9rETlMTPTDrboN/xKibA3Kga83sGQu/WxKM6QxJT
g+JBHdzVVQL2OzHNk7Rp+dC6Y2qyuJPCDs5mnQ2A8aIUs+9mGDiIfjO+Ov/mkilqm/SLyAWPniPj
b7jA/ozRWrj/9k+AXktBQSg+rgl0sif0dhLVx/hyehG/7FxfpWvzIhb5tR0LiwJGQ+vO90FiHy96
wfa6/QTADZH343VYjZdyW8ITgXSPe4RmygaO7GwUzGcR1N2jcXtHiGQ8eSVyCv7GHAxS3cmC/80P
GSSeDZXbNcxbkE1E5dQfg4qtXxWayFpqqxW0ceTZ2ohBRSDyxk3Gxtx1MmtrOlnitQy1Np/T+dM7
x3i5CMkg1U7kmFax0whWHXBjKjeAvoA4gTGbWnhJljAfJbiBK6qBEL5Iu2fFG7fBBQ/idwxVPjMS
IButecKjZwzEM3Os7UeRf7ZfRWGQm5n1HjCOUvZTLQuo/YDa3fW6kZSR+0TfJl6cq0muYqtDyLF1
P5MYY1QxLq4gD612LmF25UE1krtzfV8vK258odlLHS4Mo3LgaF2YyOMyeKHJTBL/yjhZqs2Nxsyp
h8YPr60cTxE2IvU4j05NpXAkhXkKD66BS2kfflHxRo6Y3crAf9AxDSRwg45cvi4DqxNCkEYlwce+
HxDZD+AX6dq9SMsiro905fDPGG8hxRbXPE0oHu0AMXvrnnWWKvRRTqW7eb9AgPicCsOn3RMAjq7A
obkSAAoZ108EDYqBTM9M6FQUyxfSddwQmK9iy6M8ulfTqhiEzJR1h0pjaB8aTZCOGqgra+1e30kG
79uWKFopG8QGoss2pJ0CMzUU2HgGtrfEgfJYckPOZjCDNlXun5RcPknqy2ePU6Rn1/BT/UTJlS52
tBfPFaOwovVR8fm5sBERJgxQNVIqaajJyd+gko6F1OT2KstIft6udwl8eRdfAMIZyj9ShirvGzoe
InX3OA050OrucPkUWtkstbJykOK2Qs8t7OOHrGY76O3tlptbBzzHzyI+rZ7iV1TyC52k76hGEJG9
3DDXZp8rsavOcULAWDAHCFt1l5lkbZ0GxO2jZ/9lyaRxRG1aK42SgfXcjmInieR5Y+u2VuuPGTFK
ks0faZ/pVO/bUVrConDrHfLPifi+DYIa2cYL+YmxY3fHcLRra7Ypcy06JpBcfFBd9bgggcILL1zY
h/N1g3cRYwBgaf9tD0VeSZhINY/gdsr9ExHJdrU5CHQC6d+BnIdNCJKfL/Xsvq/5ezOXO3r2XbjN
ZcFo3WY3Bv+JsuTMLYS+TCrlDAUM0mLAL4ivXC5SEeBVsphtCA5+WMKJws2N7TNRmUlbFSnDfd5I
MGkSnoyA5aj0cCTDTUKWya7tXmI2rc+0+rzl0rg6geDEmni+hnwHzkLyMh67N88ghWi8KqNcBI24
2lBtY+kVJDTn0pYldeIjGlV+5Ds6eg1zTFcl6TKJo7IfdRC1jU9/tQIrcg9EGyLInjWeyXIZSam2
YUXD8T9P5TdN/7ODpIaymB07W85+Aci6DDPzLxBthafMqq0s/xzbjRXReY28fqWMlhTWtl92Rf3C
92gSt4sE38v2zNrxbX1vtQgFaz8ZNM/zJK0hxtcZiuoILQAji4NUtlvpg9pW4B8Rq5zxOE7t4XW7
hJOAS80eYHfMJrXy9JO7+KfqYVQiMcvSrMXpOH1bwuhmScgZphGkqM6w5WlYJAt6lngSs6LDvhZf
U/uMSaW2whDBkpQcT+NX9lkrZ6wOlrjDzj6TlqdlmK4lYql9Ys2GRA2kstvH+nLp21hZLEzG3kIl
XKFemE7OAZtGANBjlkrrIzOybtNCIQOccGOEkolTnywg4Bj/rdEB/DHk1eTYZHhdM7kPMWLflC01
wrfrmsEyE6G6f/Q8p1QN07zaa3A8pzt5NC89thDvyMNipbiNLilVTnvkvZVpekMAMfN9MB8Qg/nu
QNb6ltTOU3vMNtn2CQJ5WoIuupvaHf8Wn8ar9J8aM+UEYK7WnRSPkDMKrvEqXMpcQ9IqAzflaocQ
cG/VSz6n+CfKXA5QzHM0+ax/unQrQy3EvLlQPKRe/cx13c8pcTQK4cQZQwX3wuK1XiaDwjaywEbn
bVI9+opVPYn83oAPp/vsfww2QGSK6SlpPaR9m1NCpH0gPF3Zx7i2UeWdmzrCHA49GDxLAYD4hBnb
DxixT6rAhgJm1iuAeLVLzo9UVqWJP6YUKJWwsienKSo0qQ66AuA/4mBca38ZjQGPUDUjPBAHyDPU
aTh6V0HBnZ1xir1GD9flb+33Aq7eIkPqOwTx9APKEqNLoxgHno0Yz2Op/w6siQZcMYPNIc2DQVFl
B2saTKoA1DjKnQuuuNtJeS1etPQkI3MaUCmLnNnODe0rd5QdfS4PCktNlaekMLjNkmYxeMv5y/B7
L077bw7bub3gqufOXV3BfL6vlyhBklotNUn3jpzi2/IJkwzOcYMA43lzJPLN87LiDVN2+c9GgLgV
y1Abfwq5g+PDMjOjlvDwywe96vtdkLy/Toi9Q+dTCl8XaI085g0SB58cgUOyy7AKn5mmidqcYnSs
7f/Fe0b2VJ9X7zZYYEF8kSVmQQKPorYTiWAkHentYstqnpoPP0zmrq40T+3q6NU+PMZkAs7E9ihL
CXWyVcfMCuOIt50+aLWHBaf7ikRR7VNvoRUW7y1l3wfExdXf/YN8j3H2ATFHJxi34iEjTfBTMVCL
DRdM+vy1e6sie68/IQjBF9OYsii6HSRJaj14h25oJKPc1a6C9ERU8OUNCvcAj05gRQqQNQzHH2Eq
dcD+vxMu+VhfQokeXzuAi1kAFZQZchKLp0dnfUeYumb/F+D3SkkdtHC/0SrNvS/wAbGtc7nU7uXp
OGxx6dtx91XbM+gtEpLCXDmE62GnjhNio8SKPfReFyw3jparJ/yHT61vbwjn3/BILgftwf/l/zqx
KybBX4Nrmgcs37GJPPAmLWVWg1YiXMQAFPZLXw27vfEU858k2/N7LdE4z2W1HhoIizBWSVfad5do
V4kGTwhaHBpSGflNUrlFCUqjgjGl2JkBrjcdTTAiQSkYoJ8fhVWMejEkw2pZsbqq3nIGqLaZzwFw
mlLH3xtUb8smlW8+yNBoaDPH8TXRD/hLSB7gs9Z17MI65MfWpx2hxLiAx47n3snFoKc7zQ/SR3PL
/yFzwHWUZywj/aKZoOrv2Og6Oto/24iEp+g8VUwWDYvy7Kh9V3hz5hSAE6F8E41xbzlnX6mbdL1s
cxU9QbynVSlfiPtRr7/41heoNV6VO6kOFB0YDvqz6Bzv0s9VfLgQt0yb1rhjIN+peQAjQ8m/wRnm
1oqoR0w3DSY9AjmtLW87JIerapVjQo9JSARe44r/7U1h2vVk9i8yAxa/XraGu6LUYxD1j1p1ABaa
Go1dCpRnGGGicPSdlvMfF5qdroWHA3AMzTXzHRvnFiJgJtfDaS919fkfIFbQWDY2/alYZ4M8Po/y
l2L9ZeMQJotCw2rboUKGFN84fZI/Bu1jNLEzjv0iVTKdbJJXBQiJ6oN9Yea/Ei0lS+R5MC95ie6y
0TIVSsuB4LChBooUf/AX44UGP/SIrGtrKnYtNMHL/6vqtaeP9W44K0CHgI6J97Wp58L2eOS4Hx8N
jWcMnTBV4+FQIvOapVTQkoXFPa0Cmvoz8aUty2rQtGQfEaApRydO6cDl96UQmVuYkoMGszXLiQLm
5x16JT6JXZ6bqApJsCfv/otPP7RxLhaaH93knvb/2AL+nLjA69P9WLkm0+lhB2PktU88PgJlAAIb
tX/f3c5PRF/u5SixuFIXBoODKfjFLPq2N5yX3ElP7AH0yrB5VMt3M0955iHRMWzqq3fNK3cOGO1U
0qiyXkw3wAzQUOjE0XvDlb7lkRjmthz3MKN4mn3BUCB9daWne5O7qRxPBi9eixUqoYvyoVtruhby
hymrKn8E/3YNfvD3cP3TyYlYVAGCvsH5DydM61Vyu7vFGdXsFp+eSZ9sglhpo4gmroKAZa+48fQG
8F9O1TMewECImAbivJFYld9vBZpEtpp4ufnmQGt7Q52WmZmRo5M+5nT4IKUOkWjFQF1ZjKiOzvpw
OWMC1vlV9zG3cZh1A14LLYb2U+pgFD7MEgUtjNlLanz+oWwvPAQxWyX/k4cq9Z4ALqUHMxy0F4gJ
AIGDaa3t3ECKkFyOEvXbhqYQsEkntcOwrCZ01KiRlyX7h0SjOA4lVy1W6G2K8vvndqYHeeMV7/Ep
2lVVZHK0oG1Wd8CyNjjs66A3iz+3EVgCfwNphcvi15kgdwHU4TpWG6e6ehNqXY0L2zyhERvIJGy3
OyXQrq35lwBm5vYfenYv1Dal0vLXPwUnsRYz+dAb23n9uRrNPCmrsrGIyeyQNJMB1+rncVEYpQkr
dx4ShfTUI+N6qpiq9le0KhnyFK3xCJLw2miz+L1bn3P8YTC8CRYLufasUq0MGWaY9uq0kLmRX7mz
Ih6JygkhQGKSg910AFEYOofn2adtvhm/e22yUxt3jO7lLbZFtsN7RpE5H04COGGX3tdokX+YYv70
BdWndnif0/NkOUvl/6J+rgX+Qo9ROM1pHsr9vRtT2hZEnRWAiVIAZPwcRaB8qB7a9DdkcSwQ4QzO
mCbgrQY4wuq5bfbR5tmrjFeNLaFLsbu+fZ4mwIOdPdsoz/ncFp9F5HzzLTEFJus6OWqjK6BUjpzD
EsBxMuPS8plQcWptzd0mG0eMsN9LrMXNLZsf8Vk3ZXDwwMQFjUn+RuSluGllEaDZfyg/C0pMeNC3
ha2dRByBNMpM70+M3kEOBRSb5JXySzduSC+a0KD3xebmz4vdZxLUMfs2KnkWuUItFb8Xt18tB5e7
LUMhsrZSTCf6x3tcy/1xIaS/RVVUdEpCy3pP/QrxISS+ItwVpkXcwPepbuX5jLn2OGcRvkVXqvML
1f8qie7BKqwbPo7B8ffHJITzATubJXYkmYV28qg1KOxURNmx65D7g6Vnx9IwgZ336+W4ui5bemlP
fS7okXMr6XzrIBjypggD2RS2AwUdl3E8tWykogfYjm8plU3Gn+E+slOUFB6gSMqjB436bPKIBB7U
NkYVTQod9FhPVPHuufDTs4wZEqOsBuqhPvHcJ4stNpYLr5Xh3YsJ2fLZqsoMg80QImqjAyKysXmF
65R89/hnpP657Ji0fj6A6/YpVPFkuO0V7dTSH+ApcXoq4zXBQuQLOM24KjDcrN3TfQaTufdA8Xkc
h8HZjYmsYMuMEMbQA391o9ssYVrYAY5MxoFvUdrBALfqISRxDa1D7V1e3oYAR1XUQEXa/EV8EUIJ
iS7z7BmJ1xxrHC6qoNit4TwQIojfXRB0mBwq1X0RXUxx8q1/9A699lUwxHfk3EHkd2X264SOX7J/
i9mEyZ5I15KkAa8zbMQvG9eKGMsaW+M6Q4WYZPbhQRlVuxaRUppRbyX0d6B/unE58UwU+Fn+k+mv
2YvK5IgXmiobW0bpft2j5mKuJFFUtYRJ3lbRfzsR758AmrYpOz9GO+WnIYkrAa+z/QVMzg7n9UqD
gxiajM48dHoTEO8TKwZX1I6t7bTIr3UR3yWQMiSutKOX190ACprWV2cc64HsqL+brkOQ6lrcrx8G
guogXcB/m82sA2hHlbpUURE2PvfncGjY3GB4B/DI+u8bU85BvF9Gm4oF21CsFiyPzJ3Pg2VauQ5Y
xcvu4qEiExYuUVeg8r0XeXoDW/HaKILQqo8ELhWjRt0N7jSvht6O+h96PBC5IKcgbZWwVz2Ioxnh
v2oSAWgnfpWJZmg36JwR/XLkx617RCbMg09RyO9b0TH7Aa8tU2MS55Khl3fLIvl5xPc5HYePzdfa
r1M5sEUAfIh/aeAliI3EwCCw5kLkn6ChnF6vtl3WrqHqufnZ4MjaUgiu9OtOitL+VjGbzt+iGeAU
ornRfHTrxru30m1eqyyxZV0657K6jLIiBmlTn+0AQfVFmFbrUd/eZy23eWuE2XvK18+8owiztlE5
0PCbpeAC8tWMz/qo1MJj7EUHZJNM4PgOYF/s0O8SisrRAh28WqwWmNj4SCaZ7feMpIAdzngGqNWw
cJ0rSso5ZkESjmdpB9TvMv/7kgipQe03/m/x02obQHC9th9/KaT/EWLAhr2MM6io+ZYUdZwsEupv
Lc0fhM+GU49a9Zo+a4iO+IxltHI0FSnjSem9w/4h+iyUeVs6pT9UaZL2VeTtmldRBqygLci8tdNK
f04WjVTwFo2hgVY2Q8bLi5eSUZF68JEmcYUX6meKpqP+eQMDDuZ6q6T5JbytNDuB27qXUcSirLJj
h8bfxSbrxNnSUfHes8RjyCB9Dp2ZO3PViddsoYXEvR5AXacWg3I1pfqYVIiier+Aanob0tzSaYuy
AxX3wc9X6p3U98bTTuibcVOBVt4QL9UoCSjYZLeuzVzbh3A7kJqFUnPZ1czw/XahtDPaHfK+Pn2g
qWdpwcZbqbB2oxPcxajVLG4hIOVe/4SHw0Uuh1W8oe2GSO1JFJDAPmnz3tQa2u4cxrQlOb+jwfqo
nAqALX5stuxUzg1bDeZ76syXAQ8ZhWTlYGCRB5L8FiwflMh8R6PZWvFH0YPmg1pyOfEpkQUND8Qm
poSzLAg+NBAQmojxNKWSxI3KjwjskmJY340FFlIFtYKEJQXZZhiHoKHh4D8ti+inEmQMH5wMV0hV
8LA/UTKy60pE71WVxsokqbdTWW4FZWC52S5KSra2syOwiglvGhB4XuPGFo1HkID8YQKbVu3giPM9
ZfEESwIDaMsamfpaXdMtA4OhdLEk+PYbelfH2Ftwtbh0s1HOxstc8BZhOHXWAqsjc/DWx7Ka4QGx
b5bSW+zj9AR+We0gW0U90CMst1glKl9MbYf7ofNrPExcn9ChPVJBQI4te1r37+26a4aamh7xsDNR
wilCrlLj72vsTVmiKGRuRQ+7MbtNKxb2ofHmFHbwC4idSH99fY+RXC2aWLHAzyNyf++LpG1QE5RK
W6SQs6Z9jYtxo++ozgXOVNIp+L1khoth5RtkcaM7v7MG91Gisp5LYCT2g1E0DKfMV0VuE4Cs9t1z
4QVee/SVlH7/zD1yvSbP5xdmBzrCtIvJn+OlBbEqGm8qn4E/g0813cqXeLrHV5CYePYyKctmoHu5
4wKZKFGTROX2NKVeKoUMfIvEZ0jqc0GoRMnG+WdOr08re69aQGs0H9UV9IyWwmatIOOqlrcixvvS
yMB0iY4vfWDt+Rm3bnYHxUMXqOj+nbSoOZAkGuZlCKrPliNNJMVZGG5CP8jLSUD1q5dGuWunCfPx
Asn0vUCA8iI+U4bLveIKXx1SAB2lhkpcaUCflGAtBN6G7S/xM+O8lTAwYrJudKLIzjy087FlL9Wp
7ASnvU9h4TTGOcPGZN92v7GRuRzDJ/G9oNN2dctEUl+acdHHqKk2FBCXQFykqqJm96Zay//DL20Z
NuXSJ9hsXn0C+VyUbRdF8vyuO+ze9bO96xd2nb+EWA8wCdSpepTfHS/9kGVmUzPm+fsQPEnlw3sP
H4/8hMal5RsQFEREkLGGhrtSwgOjroSMRMgTTVPdFVSd8lxPSmGH1HBV1p0lvjAjkmusjDiayrPL
rnf5NfiYemvNJl/PlZJ37T+pnFlhpJ0LqAepn6C+gyOcVOJLYGzpcriQMLzkLcUAfyLbZG2wLtpH
wDmDNeob2jqqu0tQIF8VL8U87w5HXVj3MDtPOfaLBuSZONM5aLEoCS0cvB8aeTEkkvhj4++RfBTh
4SG+kXWgJlPrgvgQRIpm1G7CYWntAbp8cp6YF2mRH3W6X6qKfTRKW68HOCce87VAo/+BjI5PGdZp
sTcMjN5RcEZ8fZwiwPnbixPs3ShtxXbMIsQeXQL/IpAiiItMhO/q1VzE4SnqAokjXXXqUBkgazQZ
v38xi7RHeXsNkLmLkBXljDw4FFuYuBKBhUgNZmti5LEzdEz2GVCrwwvT9A2hKO9uueqSgbJ10yYy
3IBnpvjGpZzAIBVwLJu+n0gtF0tASFgEk0FJeUG7YBgFFwUxttvsE5y3P3i/PBJ/LsN448utGYHL
vMxixtFShQkw64CWgNFIxwqajs8bUm/Rv1vX57t+CqhCwvZSNibfTF/xpAWG3U5OZLhXu1yFaeSx
zu+LZXazrBWl25LTDpYJZDeswWWXzdUX2MzisPCh2I4izMBlgjCAfDHUal4G2yqMZhyQqfuBPb7l
s9PspPUAAAi7eMNMd8X1bUttdHI9RDw+POdJzuexVwbd7BeTMZ8rGovmrGE+pQrUh/vztmEDVcKH
198TBm/c2KNL1lkDkFqiZAD8r+3OnW15/bxHj3LFUEYnDy2AdxGCBUXKvMZWXw7zpFLC/g5CGbgg
j4F/1RJgIPZkouWhAzcAXEEE0Ju8F7HIwPpXSS8nzCqTYysb3QhUhY6O4vuyKAElpNXVZ2rpXqgc
8vRF+/xfjYOR28o90LKOgrDTT3uCDhXokGCiU1NItKLKTZVy3UYMAucUwYGKXBuKZ/ab0jrYqXWR
aRfaTjrB5wpzngngNyy/DzdpPbSi893WN6JZ/S1DkWoV7z3OSKUQB1IQ4gZ8zcDZ7iZ6y00crxQ1
nuYZNEJgJJUAYohnAq6tcdkE29pK/kxxJ4aOUZs+6MiBYHGb/nHF5XSN2CHs78RTypBkBpMVfKir
jJ11oWfvsx5PLFkz9DJvJSS0yWH+dktrMO6IpJ8rQk2MIyxhklMX69l3sbrcosWp6W+fojh1xLA6
0JBa9TDITjs06MfIivd+G3hlmDhmNAg09Pxrheed19h7kRG/HuSTebep8VFSZDqmB3E1YhGOw4bd
oJAkmnNn7ZPi91Mcqo3+3QKgfhlprzpi6E9COxJzQUEk1PPQbFlveFGKYJoMXD4ijBIMpVcHkvsa
KbotkynsKT9NaEYDcN0hQZQiTifVMerjNCxHeAZX8u4Su4jmGC0H+hLgbqhunLqbHetSo2Agfhrg
HMB71WK74oGw14+743NmpIEV8Q9nn0LonPk88+YAnD7lVNlfuOndpNDzFQ5dDKkbTIWqwGS4/hUT
zHrJ/9cCvX5GE2Vpz0Q4mKBi7PQF+8tv3g13JMsI6c7J72Gzv8EgCGK8D8vdB4Nmor3V4gTlxrfc
bJR3QcO5rw9tGdwlxx+lFkPnI/oCIriE2ibOQnLXqWh3eng061IyOCowCmadZn/m3kGDtMsBU824
M/mh7N9PiUe98Pf2j1i+r0AoiOuYVlF3/iAOxwLTZAWFMa5pQ3zEqNki7yi3moN3MijMY5rCurzF
2+tL3vGRSlinfPLrHnkVm9K3Py2YSHJ36w22nEZEz6DRahUrfAt0s/FihkJq1C7WEdi3eSHV9Uqa
tclgMvQgAP4rdjtFx5pQy8rN4+o7cy8KwN0WBqBl8K4WIwxS6HhXNbUo+dFTjgqqAcl8Cyz7ENzu
N8QywVFsQuTrglyDIKnJO15yny4o1Zv77I8GWZ+KwXz3Xsth4pOTtnV67cwVNHDRwaCwFCaOK9ld
Lm+1w821Sc3F3gKqWl6vHSlCRMMIkOrxPj91QJP5Qo2do5+G/KxqdpEv2s3/1sYZ8ck8JnkEZyP4
61qoraJOOA31cA/tK/XmGQkL1LHNc2gbVvAFS89lB79LZNwQRuLYM0mO6a2n1Mywc+cjEVlFrAMx
HaIlqAXLgjGx3POYG73SOBb/3bdGhhxithEmWK/jIha2C1gR4mqsBdLMUoE71vCmHVga7AjiRisq
W1MW546RgVfq/hyBQIBpJbmRAdGtd1tmZm3/HDV+eRMmMcEhPHYDr+qe2SFjF64ein2e6CGz8hKl
O1GgQOlLDGSvLAU0sx05C5Fe686TxPMWJYk9b4K/AfYUdKrd3ogKhYKUQOV0JPXO8wY9p8GpNlB9
rzEdvsmW8DUhCXDzLhNfcS+GdXqMcYi08cr/8e/Q6xX04QlImNrk46u4bvxuDDQGl/tgpiX0imsJ
sfeoRJyKKc8cU9vV2GkHbxXBgQ0wbDaa228Rn35lzqGywIbky/XhI2bEA8e6Jpef3gHu6mmJn48k
5lwOje0qyX9oxqs9rPMKDaqoMMYeBvyDKrRhMUZBeu63gz0+Y3z1l70hnmi10KsBUl0FTjjOZluP
2sLdg5HaOoum25WTassn0EejcWQ/2A3KD87gGlWavY2DFpJzwBx6+euJSGR5YeajkrQdsJuFNDmi
RlZfNx1yjJ1BdPXrYTOOuBPWaRzfjK0N7qSqqrI+lQ+9T3riRLBLHYUB0fg4czFdtn37upxnZjvU
qKb6A/ONxxFkKrQDb0n2Gen7lYkLdQWJ2XTUSy2GTyt4Kdlk/qwWKxHoO4FcC3glbgJ/jl+fpDk9
W7OSoxXm4BcLltQa7YI25LYcM6fTe531Oa7bnivzM51qMSblyMhYn4k8jIG4iBHh16gN91/1dALZ
ayDEDQke+EgegKBmuU+eEysn7WQGhh16QAYYFDLsM2vCVVROBNApokntvL2T4FQhPO67D/tTK1UN
7NupCRI/gc3G3Y0mmNmB7LaKKAUTcT8ks/43j3ybC4LL8Ewe6cs2T4EpT/s+IN2n3+7lYbdAvnnr
XEdLGEXemmf8kzHA7X9BDffByo4hBHf+hA1Wz7qeAfqV5BjDNBnBE4CfeNjKPWXQtZ0DG+QNoaOF
ZtfB+JTbL8FKkNtegmWHhstj9QokhthgcXieqp+d2HmQ4oI/7YNGNc/+9p3iCTH3WN12zSlqCM1L
VxQwzi7mtBLNDm1pHidM956vUn+K3SbKdPfzsbiXAVlZcCUYm4R/gMNtLXgqQWBbbf9H0WGIwP1g
WTQm1BUvTOpe2wtFDX239j6OGb8YQJEw1/YvYeodECgZknL8ixBFhd996VcMnpdq4dcwlq3KF5IN
KI4kkoJKVmpFXAf5I2ZWZgnSCuw8KVpX9ieiwi1FgUwbQVAY3o6srJKpYIKcqreX2ERTnV+uhiM0
1w5cZfYgTZoC/9VGSC4TLh65OQai7xCvsOA1dub2hr0ahzNLdil2LtdNINKSEOX9fweHg4kHQaHT
iZvBE1afXQYjWBreC/geacmu3byGOQ6TnX/3T5diEuPuYE1cHRdaY75smoCt9Epv40AAXzEgqwEz
0bSbrblQFztFgVuTL1yWHmf24vXjPvb7uROWBKEVxriB3YJWGsXaJ3zGTGzVw8jsKChs6SbQK6Ov
iYCPFuEqfJya6n1GUEFkOD/nkv4mm0pORUgxFoDz0YpnjmYEiLdUPNMpkkljTPK2CVpcgHilEu52
jlYsCyEnj9fNgYOZXi0i2hyKxWKEQQXecbiJUQ/NBia0VQPm8gYWl6DIGA08t1z6RtcWANGQ+X2+
MUcwluwkernZcUWm8FC2pW28zJfCwsGSmAYwSXZ7jP67rMRxnOYL2y3gpKKvNhHV7zCi5/QunN4L
P0qFpXFTaLI3La3gw78bDSNJseRQX/GeiFD5On5hIYxAQ3Yz2zFLpfN9g/ulwZ0aa3C7yh5w4jsn
qZ4z4kJiHeJOm3DrXIITxOK1U9+YVX7OWEv2kxvp5RCXJOebQiQEySrQItjueGouw5/WKmgf7rLo
iOWJQ7jSiNeKJIIK9RMir1KBSP9fsCt16XibBZKVsOdhqA+tdvS78oUgRxRbwcdrvFfUqJqNdAk3
pDxJlc0hU/XfhYLUCQgYwDQKN4l4h8JZjIW2lee6k6fB9spHXcicEWcGVE4QCYd6RcXUQINAog3v
xKbaLTlGuSttCsHWbNg3h+olSNqJtNOD+Ew1Ah1Dm6XOJ4VOZOhNwBBu4NOVmJ5v6iuwqg2o9Hbo
j3Rxrl/ZQcDptlHPx5DLkW7O4/YNw/6HtxEqSYSLuEGD1BYB7w/AJtYoFFKk2gb1aAeUveaPJLB9
DgxHeMNRESAEE2OCX5QpaML2VEf8pd/RCEOlgfjF4YEvXLitZX7TM7bzxMLmNTp4Wv4d4gKrU2K/
rI0XivBvONLCdElR/3Z9ZOo/GV2vZS0BrAsq5WtB0ECc+vfU+DleQOjhxtu/3ZaZfNVmBl+iQZc1
lyGMRqeX7aFS3s5Lwi9lKQ4rv5Y+pYeGw3HG0xh75Yd9mUxdcxzDzguYeTwsOaPvPKP5f0Do1yHe
ORBiYfOR3w7ucIVj1/DIut4MivYcNqpp50QQ3ZzfCP1R0p1DdjLgEtvQudLe2CKYjGX4WOVNYiqS
5yQ+jrLhYDImH/Dd5WZHYnC+nR/VvqifRyqc36zbSz1tiqUgXFNJeCSk2VB3RGXQvnQJZL1V3Qfc
qI8sIeCAb/wpizYIYvTGcyj4abvZ99dxKZkB4dEbIc214+OHcRKClS7cy7QCYt4JDB+ossKCMYMN
aKrZ0JlKuacBqL12pNziQSwex4fCZz1RgFu42upcU+4otXrkLkcMsxhAjd11GGYn05MQJD7cFg7J
KKoaldzneBg+QlsKriVBGWZupU8E2yrBRePT8KgML2d7XTrbi/v9p4ZoAQNIYoO+SJRNmKbYrLIU
c9WfoSljJOwo5OYVEf2yXYTfn5ZHUTPOjf3fkgBByR2gNQtDFwX3zzGnEBFYqVdMzyze0tNzlJB1
si+lpIkXUemy/uQ5cMgU/ygOYrgnth0btcNNF3sNty0jMIiZRCkG9LWh2VwctXwxcvWRxg1K6MtB
/xk6zsXTnDnIsKaD9IIP0NbkLU+0tFRBxsb/8SWC6RjU4M/fMDFq4faDPd6yPT2PU1cs0vjLnhiw
4JlUtAU2y+p5/2RRXBYHS/AFGGmkhComOzQ605CVRbGDoNTvc/H4Y3Pd1hsAvl9Kg+9xUT2+unlv
9ZHoVGWjTm+tW4PZmV4r3+ZhzGlKsAHUahFnT38yPWHqGExRsik1ux/trbjmvbodJVBG6P1CblqZ
K8Zt2Ibb014QifqT/Wb9ezLQwEoyXzFvvsx6ht4al2LAiofcktNyuxhB81nyNubJn6ojbRo/yEDl
AUqnuMwU7qIDw6W6gnGJG5UC1LcXCfe0/4+boUMPqa2Aw4DvIBboJEFCcy5nddu5FDBVn6w3Qxon
DCuf71HE6ByNDvsIg6ur7hdyNDWsAYbVm2Ja53tgvFA0i0PbL7yh7BT/Aa5h/T5OjVucezd318KS
lNak9/HVNyQQ6YuPJq7tkkzGysG/S7akW0B8FTe3J5Dgt45eCP47c7MV4Zu1rpJv9kSYdFo02+Qf
Cvf6Gee5GVWkmIZFpgMq5W7nPm3Bjeppu+HKumRDmy8UFs+qVlNgFbRU4pUowhLvNXLpt5aBJJza
5g7eL1erRDwRh7Jtsci3/sZl+TYXC5kwqeZGy6qVFr1cGq3haPHtHtjo+qXo4GWHFS6rXTq7Kd3w
X+45WHZcBgtHtDBPznVK6m1KliC0idx5pJUw6finHw0aYyDCTyL3lXgsV7OF0guNM+pvAF0NaDqy
6eI0weSW9nTR1psVeDfvVeWXA8rSWIEIW48Yl8KGkki0OWtgH9zMpqQ5Xx6iIo3FiRwSsVkBYccu
rIM48uVL++l6rQED9BMfL1XFZDIXXZkn4ke6V5TifTPH4V3MmWkJhkaoMioY3PB8HILYMhwHCkmf
9DrzZZcuxq+GISCSLgGr8z+IGNWaGqthl7ewdpF0Fbnnb3Dp8PALuSnY/hHwjJkJcaDiwNfVYanX
zj4LZtPBTPE8o6H+WO6j1sOvK+KyTn9P2DPTHtdf46QD0Eh66W6UtT7xTb8mgJG0efJqzX9oRMlH
u5fV0qwb07gZCUoZ3TM87tyQpgoIwBoKLxtj8a+rF7mXvocNZ9bUVwaSJ9G5GrHL9YUAnuHoR8VV
rPfbsWv8Hh/vsb2ZriP/gPQ7KQk728RBvqeQB/FartDSVC7oceQ8lxgcTdchfq1nQQrIrl7mQn3W
OPfWf2vm6v+9fKlolc4ollbVGBROD5cBKF2PkhLg3Km75GZZwHry/D4IS3R6QVoHowBFu9LCK8q4
uhisOW3S1/CHjAf8dgexHGZhiQESY9JycETTDEaIOgx+aJuXIxzRYTLdTw9UMtVBAlUQB7+LMabM
uxC9Mzrf2bSnGXVmSTbWLEW7ic696YZkBjXGEt3tKoCHdUcPAXRgbHLo7Rp+sFmdVV5BPYB9qtzq
+U9Rfy+IWP6FCnRJQdnidERy9X/d0cmYKLDPCBqCQNNpglgGF/xgIC2NkdkdfIUh8ORW1he+6hw9
7VLpXfd3QD8xETY+XXLGV/A+CaaAyGh4uJ8+sARXZkDRQAjS+688ruBsu6gRj3EQabLYVsO0DSxO
H5oNx8y4BeYm7SAyCba4Qcj9S1pcK1q96cykC+9f+4+GPmyVbKyS3XGrpmFyOVMha5xEij6Hmzov
b833qU57TTgKZMXkk+GJJxBrQNj0edSktmmAJGhHtcMy/r/cVvJSRwnUmZk6b6MhLUhXtfkcpjsL
aoj3FuXoXTReoLuMkY3hgvr7uBkk7Nb2XcQgM3xxdz3DXxCWVMc6iHlc1OAQr0eU2rkyfg7BCLjg
KZLQAW06/lfZ5CP1LWbT2SRdD5hL1RBpMeuM4wOfI/169grIqsVPv0oPPGMmJdgcWkcV7FwrFkd9
y7TL1FLAiAp/CEHr3FVNHKu2A/n/2YHOrSbavoWs7LESHUoxZ3SoTrvA5KJQecY9K/gRLW3jFZJv
S+2CBmDpNgnUqsUcQ00bXxaaJ40nFTjWCanQK3FOXu/bTbJyq71O7YpShiyEok4fUqCVooqhLXr1
TrOeDLSN5H0gRKqz2j5dWXt3srbNEQk3oDvzNyj983sHvC6k4eJQPcBxoq+Lpr2mXF4YbDUb4fQA
LMK//FbbarUGAvlyYab+/TrcAPHcbeg77gshW7lZf7xtX7JUlxKiymKt68cHwB1E/nlYScK8BjPk
cfJOMaFp/Rl/RyDzpBQm5LHGH9cCpVyM4LLMtSrvcGLUI7kNeWazM2w6rrkN9VneTA5NR6f1L6Uq
quN2rxTKyJRlMultopoaiYNLHhuVWiQmYSptbwvATRSkmC3R7F+ozWabnJHB/jJABc5gMSZqCCDC
mGupEXzO2Oc6o5wfkGCyIoPwbO/bP/GgWySdOJTqKnzqhwIYjzZ3nGnRIQLtdC26TEIZAa4KY2U7
RSN9PkTv28zmTNLow9B7wfay5kcNvgwd6WjmpwPYdeTR2y6zmGiT9nXhXZIHm8b0Q3akxSzfVfw1
knpC6YyauiufdR5iAY8s7MXphupDX1L8qLv7doItDMXfKPLR4mMwpggh7E9IUCVXhAomG+OGhBmV
au6AmTFTO02/HavbY6XYtXoQgzy9dSYwnDCAXD4lghCGcZfX6u+485FkoOesdDmHxqrFQQMu0VN2
fu8/g29GXAk0ty+K9x6hOLXxWPs7YYTsjxtVWlIzX646XhfD4XRjGC8EOwA/VwzR2sQZ4YiBEVYj
dtb4yl98rc1/MVqDvpL/Gn0gkYvWE0oo+eMWb9cDee9U5/g28sDCTLIT5GOEWLZJjwN33jz0FjeK
jeQZ4Vwa8aIB2uN/CJ8ckd91VNi9xMbqqBjv1xTybgR8jHxu+0OPpo08S7xw4YIBWfYbEKnf/DiU
K4+hs3DjzonIn66X6ycjbfE3meUI2QalVJHVLOYdcL1B46f6Iu45ZoDWZOhiknCU8o8+djBsppqa
1aanis2zqcfKUWkrEr/MXUvwYmzbLc4Zi+6xoRaTerAXamNGosp9WDpHBIxfkGOUENopISd9ERsa
fLPbwGVM9HH1i3qhHF0LykpdvBMtFLY2zzw55zcVOH3Z0x/QnSg8OYf7zMiYy3z7DlVha29UgBmp
hbDNeMXaeNesVxDO5lzleitIaB+yRZMdBHvVJw71Wr91G5V9P5V3qiOEb6iPk/v95wIYf08+KRC0
Y5O8tJV/dHSvzE3rTK1lBZRAEz66ajyrC2TH+kaxwi40p3AODni1C63Swejr99j8TSZ5Bm6HxAmA
xNKsHEtb2GkOJTAp3sOoUrb5TWvI0e+ovemJLYjcHzSaMrKyONeqoOXFLlT9SfHJXBjOq5IJbDQJ
0figkv7sMvRZ3g/XHYoyEPJBU7gJUnZgjj6XVDmiTVsok2yy/hQJRiXpt6h6eKgYvUlI2xNVQil6
XLawlehHl47hgJSYoxM+hei9Wh/6hJDdh1o20hhXEtmcAbZoEH1zhq6MSDJBvayjl+816L24g5F3
qOuLgpSgy8b1kcyWDvWPyrzPZLMF1E2R6/0XU48L9ZwZ9KNDjSgs8M0HnTIdS9c7JTNXp4+oZuxP
vs8Q7QPLnuyuhlIxJb+wFNygeBk12LvHchla4NvK8aUT70JiL5rGV+JvQ4ZcwtLBubs1RCDutYvZ
PVy8WhC6+E1+lEUF5tav0opHqCPkHT0+JC1okNuUEso0G5GIlQF+nLxC9KDPa+aaFbSHLK/Iswps
pdbgcOENRLCemT7ZzKiA4Aej5YT+lpYMAq6FcclYDTEd1hnaWiWJeLXP1O3MDmVnpgRd+FjIFrPC
7Y+ef/I6VoUdsRo2PW/9srgCkY+/IAmjfGMOuQiMR36+nU3M3OQ07RS9ausN+AJMXWgzzIMUo+on
MPlcGBM8QejofqkyDZ0IDW39ri65Zq8LEcxj7lihoc2knhnLWB+ZCEQvNn444v5jSXJgLnfsLowW
i+54ke8+kC+WVxFon8Vz4D0QgexY9NZtoq5ftPfTvpknHlX44xWC+8ov7aEl7KOqPM9oCjI1OBUb
13J9Y810nFalS/b+lp4qbj+C/4kaujte9qPDcoR25W+ND8h///cWWOe2w72+Ev++GrjRll+PP6GN
lCY1fP6DZ7MCEMDsyow5pXw36v8rjj+/Wj+m68VLLhsY5zNpZL6MB+eMcoW1zA8khUjueuCqKRpG
8gtvOcrHRCW7S0o0TpTCeOu8ohj8DxiQ1/cr/uQTi3L33F3rR+jRmgl/RmNpDl9Knl4PooIDLfAd
Lgg0Em2cNvtW9zuFrd0qfvLva/1flk9/B2IgolqWgcXm9fcW2u0eJFxqO8NdTsMm5yl9KOnayA+Y
H69r5LF8jY5OpME9eOMeTzXFTK/GlKMbXBLOy2KLMjCU6h3Xxdhjb2+Gi948JdAYJ8OWFv57xyVr
2eehbjpjsM9INr5ud5OCMnua2KOoFBWS9GS953AtlrTiqSlrw5pBbvPhDJEsQM4xGzogiGGJ+dJf
2s4eSVGz8PAIGgUk2gO2kYcEaryWPEm5E4zVrIU0CkhFdqJS4Nfo+UzTM4BlPaCouMdMbHQtkGS1
j+dcZsVd1PBnx+3veRVT3xwcIHh4SbFeZzdxt/KDDQ/Et0IpqqQT0jM1LHxBXMcIAKsy86VqsDaU
mcPExdpGxxyqoghsJciPCz6K8odl+HHKEb5VAwMDYF1QZdjDKnCOYg89kgpu8HHY7MDodFB8ed4s
oUNPYqz5BXmZDCTe8RwzYCiT0eewrKYMTaowzEmGhE8ZO4CebTb5xPfAlDIJeCwqH0evDfK7vtuX
dZwAEXSPWzcnH1P256Kmf9y30NRA5dCbxiWvecB9tFIGYpOGvTDePC4G+yhCjtHnQzG3mhntaCie
hbttUWDtSLsoChrbMt3m71cs6ztlQrxefpqFEurEKb8Bj8VqUmtA9Or9+bn0W6jEz+hfh/97lSTd
MDi8ptQ296PlUPuQaN40jhayQXNHWskH0Cyz0TjgdDQxO6T1HSOyrXqrFvKeJqwoA0GO8WTNdRW2
YmNawN3KVc8oUuztRyzikVZCJP9GBxAtFdV+ySCDAbJqwGuLIVf87nGXAb1n/iMHyUcvG0pz8OBO
v2Ll6U98Jx64hvbuyiDvaaBrefbHonMaw6m82+pdJxsOuCzzoeYjO92YK7pKpNXsxKfoB/QBPbRM
8cUUt0j/r7H9bkIIgj0n+V2QIgn5pzLpY1KiBBTidtLbt0EWlxGlfOZJKJsXU0DqQwRVz6dqhCrO
dCDzJaHHl9XY5pTgfC6NcGEGolu/ipwshN2HWoscqA7b0v1e9ktkKMk+hHYlM3yiny9sYcOp5zOq
9WBb9ajE30EAnn2gdQjAxu/DNbKe5KChvTlcIBNvT1wGnsUSdu4048uCpWTFQVffBd+AAsJdDHFi
jfmQaEgLZfWuVYZqTyA7EIwk//g6JGdkfU6+HJ+T28eKByFdt9XtKCojqnj+OZvMwF/GXFCOOAn0
9mHQgqYGmHh7HREggpOKJ64+TYlPaf+j8Pq5nmQ1NnMsf1qH8FL+/ntisOjo/fgxc5JIFy8VA/EK
A+B/W7/9N5pMqrm0YIHkg/xuKCETlU48OFtY9ET2o5X2WOJ8Zj7RC0qeJvGI+xFn5Z58HKOIotMc
XoWvyXSY2b6vzhuzxqzMKBhlocuhC/faNJLLTm1NPHlCS2hX7ahEk2cIjLkFH5MbSrFXZHgjf4J8
xXmpxYH61YMbUqxpydMYd2iK4GPq2awWXAiEm94QTNntReTJmLRyfFbeaCeOTIXYiBNnbUCEqsk1
EKiYuUGME6Ex/k0YIv7VeLoQY8sePv6cs7dXybdy3EPHj/xuIknTym4sbSLEVJSc34ChQ0p0BeYJ
cDyM8Bjj2wK7+eVrk1QA3Mp/2rxwXIrbNTuRbvPwypTvic14qJiAM8pjBMYUECn0hdTIh9TMEgv8
Tq7/R7BPOJXlbzPTYXuLSR6/ay86J+5KBH6AGIBkH1Y4W3BDBk6sWC9XbXxegZ8Ate6cABbUMo/v
u+3zhI1EPewptGEnuYBW6/dePnJesudqBniPLjdNMtAexqEKdKBZR+/iM0AXjJJjdrwOvEnvNkop
tQsTUJ7UY3cgYmeUpJOqtEE3NCqpo6YCWLhQbrRNWoB/6h8tNn1rMvu1sn0viwGx1NDFksL6ZfA8
VyTwy8b+XJ5AmIIi9cY4hXKP736LSxMOYnCNz1enX9hQAvZENqbm3mIFeu3Na9pWtI8FnFO9no9G
idkkSIOUY3UR9n7IrhYmMvzNUCqAY+St+WrFA4hjOU+CunGW8R1/QqCfCgIA8JLhvDp1Ki6+cEqO
qDiRf7rLkV8TS2Dn6O7gNKD18eBq+gUaomevKYjErXh4xC/XWkGeMdxB9JicGH2YICQZxkoSOnEI
ZcXfwtT12Y1YTxZtFXZh09gOc5iOdQDK6XvF17yheouRMKZxlwqzs9axymFStvqveRFSzPDJ7iND
1dWpv4IZ28MMjeFvTx+Q5t0JpWZGHTgMcvcx1svODbWl5f1ObwuMUftW861iwQ70Jbe1I1/F8pNI
lzwmFfY4ywVaHFohniY87oTAfBrSkeGW8joVuQxdkeXP7bHNiydnAP/Fo4hI06KrwVzFlQYum7kL
vRW3zpVW54pceeC+g19KTB361YXf5Hi4pQRmBlZOXjpLkhFqd5mRAlFi1v6Gj2LeLCq+8Ceulqh6
5AMoyftexpSsZ/L91JF2SxOzBGZyiP8iK2TXjvsYef2MTZvWspFblttNCDc7LK/LQZ18wEqeR9Xd
IN4FgSBaljpcDGdMpfl0jTAx1p9gLhWqd+xK501IMOb7c/rYUaPlgP7c53enEhg6kDFbtgXndOAi
b6Dkxi5gnCSmbtYsIQ9fE9qvDjVsDdHSo0lL1VljAD0ewv66cmyY4PtmGh50bhbBWEMj4fZHUJwD
xHV6VmVHMW7KWYAyYaEvjFJVnLm+NORQe1nnjgVnQLa5RjbJZMrnK00TXdvsa3YqPnw7P8YmZwac
T0RBMawMAJQk93c5vn6kMqWEL9QbhgYUGmsJdDjRLSFm35D7MQB+H6KGppOLxTBTHJYW7tT1vY0w
opQ4mhhbBgvJw1g0MKVz+6bk/PtPj0bbYqRwrDMVQT4bpGJXFvjMKJmOgzWwnpGZj/rLe/CPidZS
VAHkeFCNJnpoZthemmdf/buM8OtpES+XOYW2ArMWVocuwoXLYlMqUjXbjLykgt0yoMBifI4E/m6P
mxQ+HzAOahp5/YjTLro+ebz3aLQRZRJDSHggc/DE6TcCHaXhvwZ6DGNEYQMT0Swu8DEP/KTEYY0x
tCxiT94BbIDkSPatH2bWdD8qB8MWovNWrY0Z0gkZwJEujdPElRPZTlS/U/ejX+Dhqheb+XAlXjlY
eTbO8kcipgQcq+PSfXns87ua7UqAs5cIjIpCMmgfPj4lhbhEe0FC7RHF6UIMuCHMT6KSwWxGXcPl
0SLXw0ZnYmSTWTn+hXOGnEms4Y8ycgvhO+owmbVekktYFn6pXOVTcjuuilWkR5mntXBuiTNt7vpm
YUaVHn3BWGtg11jFDPRkDGh/gReX3tqLReCkdy52buggfBpahV8Gf39ACNp6bmnnj7dpIC4jjOvc
qdcOshgNFos7FhAYW5HxQTjRZEP1NF4R3NwaR8Cpe34qE/E68yEzoaM5+3HAZYhWTRBhRY3BR9Z4
n6sCpMIhH/8e8EgSn43wkdZmgso9btMJ18B/UaBM1smQkDW6PL8CYUaQIW6o9olvrKaBwa+ZM3o/
jI4RI6s+b1srNgYOZu00VGWovPWtnj0PgU2ARlDk84vYFleYkMlpImo6dKlMVDhsaZG5Ri/S4T9f
JkbLvJik0c0A5T2EQhkiZOZUBsk5rpYQufN9u41+c3Ermhw7WQxg0j2f464YO2sIHm8sc7iKRn2q
UDZuBOEO1lIwpET6MoRrvc3Us7ihxmGEN/UelvdqHFeiFhaSknSrPKfrA/cvhBkQwFZPOkLY5ini
TQ/PKaFjaruinTOyeOKl21NFNIwF4DWNRiIzPxYrb5FW38s5f+MnD3v0/NULzkc4jXXq748tnQKr
G8PDOQAmj70xOH2FzMlto3+ZzvINPJdU76cDptmIB3EEWoW7holGKiPuTW4yjm8vHpf5Q6PHD/8n
4jhBX2kb39uVwkwVYB41DYYsr4R18la0OS2zZwOW4S2De3MmkcXUD9nWqLt6GLkpscJkrkuIPE5q
KJcqXYLqXktEJ8bkN9+U9hIM97xKA4R2mDiuJu9Hpr0DTOyct+oP9nwNQPiLM/D+Fg7bXzj9uWFd
vbuJYD2JNVD9joavzwTIZHF5WNd64oLrXBp2Y27piQgnA8idSOqbfjiwCahaH83AwwkAy6bAgERR
KZof0RS+JD3n73O3wdR442y+BWXjDe/dUZdBmdhtt/Z14j917Jrq4GVtZoIIbLUAcEPlPPe/2Tz8
ObdKM0E+jmfGHvtu11T6lID55G38S95zr0rK/CvZpVCkounzQKmt5JQy0A6Yx8LlQQXWnO5ETj4B
Aca0Nk/qGGsQ06v/ntC3jhkKbb8K7Hp3SJhBUanBmp4auJhoIehZGhWuKxOMvgY09XpF01VUQl8x
+iSqTkXVq3DewWx35DLutXSR6w6USIR0BlHFcR1xM9zcXhvjCviIJlzAwRgjpB8N8Kelh4r1rNpv
5gdlgLliqOjUh5FdhI/0E/mZOdKWSiIrjguroUUn+QFhVsEOkGOviNFW3Ys9DWP6Wn2yJWL4oSKh
xIgalayWqRJ3hzP2nrxc9VH2O1ghCRJ1zgglyzVVAccS8RUb8vaI/KguAxQz4xq20Tm5/OlH9LPZ
IliGb/E2B39+yO5Ntka4T8k2TQbCVuvDWQoQMrbJB32FVEvguchoZ3oRvwDPTBgeS389h5FpDPWY
nXFAXfkTG5vQxp/f6y2zqEDlL5iGuawAGKdbgBqOs/c2WXvX2njCte0d8pDnmc/5JKdFFNeMJita
plAreEq33CdMwop1B39VYoGHqx5F+XqnugzL5VB1CorxqE2o5Mm4ghGb3Fp280XLW0UxWojqV23A
pyPXgyYxn7ribd2PMnm2djlTqub3LNBL2flsv2g/8tHqN64e1zjwIQsO4My6bPr04kRtxbP83Ir0
Z5ots5hhNeUob9aH7bht9J08ZAwYUDgsQoIAApGawkMqhVgDpNrP2Gg9guaaCrmF8hvGDSy1Fcfd
l2HChojOHQFbbz+eD8I6teI89Z45Kbdws3eWKZe3b0F+85Sk4TVKu/XtCbwpPHH4RkEDvt0dWb3G
VAgaaKV/BAs04sG88axbKNIhiIGOES1Q5Gvj563fXgzfQh094csO58R92LVtzv0sQrx6yVNcUhER
JMP/byTR6+xNpT5fr4Mb5EULmtEdtRwXiHr3zwMzCMu8cqYnb6pC4OTSyJJM3D9wlLaPjuBpEA8A
TYW25TdXTG3nokeAXahQ5gChrxqC/7JIgovgJIWnUdd+yng0MDHr5v40DTvn80wWcUWtO+btiWde
yudsfjXYn0rR+iitRb/QrKZdXB4Gc2F5nJFDkaeyCyh2ELAbmDKdL3VQlLAsvij/qdp2oQdqF1sB
t7YeqKS0nBD5opYVHRUETm6tsrnsHB+1jM93QJRqn2mt6J73unx7D+QkPWAyl5I7jYPh2iFmoPbl
JeIcWRcseidVeP/pQ6Rls9utuKmYQyciZs/e+kxPlwOxNqumPzOXdSRCMffX1JTe77f4faltTuen
8eNW8o43zeDM2UPpVC+M50Ra3l5MeaRAu13UYBa1+P2xrPxI2eYfchFEsXyVoonDqFDHJ8apZKb9
plIRyYPBzjUVK0I+1ItkVj8OJSigl8Bp4+mQfMIAFWDbFRG0/KTf4UBybBhS9kBFKQ8NJFa2oqJk
/tWJOHnfSSHvgqy0Y1GACf3tMclNdx3YHZw2/KCxrsCNlRQ9zMANZJyskHxyRqYiWXD3X7CeU0/y
owKm802F5wwjRLIISSeCp/Br77Q7QRO0/rP3cxwjCuiNfV048Da4VXKqXoTBxtsdhyYYPHAZPkbi
v/4PsCSOxy4lpeGgfyUudd0yHURpLgxVYel0xijAS/j+5RXW7bJZKaJhIUPhKEib9DFDxwyGSPeq
MJdmFOm5EWnA6Mx1CmEP7OvnGxtfx0QAc8yHx+8+RXM5vHPvTPyQEwbA2KlsfDke8Vc9UK83fGNk
2wvyahqVmm9sAPoZbkRnsQ4mpBoBKKhn4kv7YO7DXXbbkX0ACkLFfWjs/XZIO9ESCfecSSpxdJ1U
2j3BhOefZHcfE3CgnVAv9wRNVk0joqF2tnDtyDbTmO5kXQisBwl72Rx0APVZno55J90hEamNNwAq
HktfBr2K24JVpw0vcL1pzKVyJACBIjwfTUhGaIPk0qKqiEVq696CIH3Gtk+EsUhDBHsviZu/HbQ8
9eK4c3EDVQ1wjcKT/ZeZxhDHZymjfnDmJI4lgFSaC4VhFeCR+l0MuPem3EpaAmdKXV9hAjn/KJVA
IZAskTJuvIKXFoAAJhM/zytkt72hA8JRa5oyYQDSwk3ETf5ty5l6E/TX9mRkk3aaUQUiN8wFEKHc
2pkiQuJMPkLTnFF7a9w64IMIu1f/ELIR2nBntaPSgAqA+6jWNhTp9fysg3Co2ISEmftuDTF8XCtK
9oyLAuq5lGoyTpw4p1DRg7PWkvQW8gXmTRi2EJ6iABRXHmeQ27kZdHYxDZWdqkIAnc+1rbHsljay
7rc1IHuIywkg232AHB+bwZ873vjIhWGLxgZdZmyGN4HNGcoo+II9WwyWSNuE/p7OIsgvI3FXnn+z
92hZhJTy6bieQ2IFo6mxaYx5zh2N6Ff7Wh4enuzAja+q//lWbHlvY2pqJALvTp63xHNRwV30vXP9
eQATpUK/a/tWsZYoJ8M2Gg1hHPL9RuNuQaj6tpHv9em4syjjoTphswlQGjl+tTwVuVICjQ0Ggq8V
GQ8dPudtDjmz8f0/EBboyOUIhzUY2GOUk4sg4cJ0U+5Kngak5jvgqaN9AMS5H1ZaI2LPPy92G7hd
/JhwLzroWLajXWOlWYCJO+9GCgogqsDPU9eoFgHdOgMLXkYa4ZeJhlX++cCqLjnD6J3T4cgoppGW
AbUrRttqQDHnscEwlI8qVisUM/0IkSMUGbr9uQiEQYEVF6fNT9PhSf4FPptC7VHRrSIwBhrQC9m8
kbv7AtHUmZXWq8HBE4lc0SCsgFdCsKcv6gTiNwdYiGQQ1RUCt7DcY8p2ePLa9dCIJzEjg5subLCK
G7Hd2c365iwGvjQdeS4QfEAqglaj5XEzA9q68UU9786PAlOJLUtodiLzLn5NTexHDGa6zbgg3++z
kJHvAkYvv0dtywgiuS52vCN5CWI45vdWkmyx1wXy+xg6jDS5sJxXapSai69Wuk+2vZrkwYAd2pba
MjARPK0lchcy5Z0Xw2QCkjYc/A27yd/4AxNrihp67UGgKstVw7vjBY3QAHjw9ccGgnC+WP48L7dZ
PTfrq4Ey9emp0T1oAVdHFnvgCgN5T5IXZlVFsoKH9LE9mQf5wFlEFrIC3ZYnGs006iXo6Rdbn7dU
q3ojH/Z2zC4cuYyXSyFSgyFjmF3L19Ltfy8Qm8ijY4OHo1NgJcTZdfSjVPZJW94ut2kEEZJzErUN
6xtuhI1+D9I/jwsr6Sg/RHfs7L+k6oB52+hbbpa3a8lJkMI4viW3mtwQNOmf49p6i28t0/nYR1Cq
qRYAupQm9GgiUP8m7Ng9aq8mkkSxc4WhsWns3Tqrz22pmSAAC98tyG+jhr/uRu9jcF/hmflrLWX/
/FGKgfFIBkhSucKNplFhIvl1+WBFpohM4boyyA6SSvhb1TsceMe157uEjRruw0CsHpjXEEjyp9r0
uoyhllCNQJ9+6X+kppX3/0NYrpjGgcH9TRLbPVCQsFatyUORTU9MlQ3JRsCQc8A7VIv/rFuieL3x
Hlvy7igypxhoofbM+0nv3TQZjHSMTgM0CZb16mi7uvsqHw6+2lg9LIXtagxGD0MYc7TgisN2ce2D
kR9Mic1PI6Qb/9Y28vQnJzh0AwEVl9uIVKs1D6KEkH+fkHUdDCbN/v2tQHdV8j0GsESVimAs7fWk
LtaY7kPqO1WECKIU9tJU9CzPcMPeK30eSjcQtB6aSGtiilADGImtaCFP4lvvhcEHnyAqO/VAI1dQ
Q8IWYFrr0M/c2dPdnyj9NzbnazTNWr5/ADzG//abClwJ3v8cD2HDVRoYaKwyTUe70/0JjUpjKdDJ
fy1lqtzcOVgmlruuMD3yHnOeLhlQog2KiLaR3ee6QDpHPGP6EU7VKbshg2r9hgbY7kNRpd0jpGkI
MpBntPiJQKWFLCq1ruJwzaoGXo30HuzPi5a/0vmTHoli8ddV5OsadvzR6O79CUyvFItCM885tvlR
Merl9c4pgOrst84g0lsamw4JF8Zml8QeaiWBoBER6CVlH16Y0cSxZCrXkGd4spFDQ2+iz+mFeQSn
C5ZsrlHXof+y8b78gVXt+hS/thY4njZDwQZhLrU7Qkd7PbWqHT86+InuET7nYP736zP8SZX8m4dL
dX0y9T5jx0obdLpz/xiaC99P9GXdAu1l8Uqkp2mEvuXFjj/G2fWLh/CLVNeKoYkzHFl6Ewfy+om3
XC9BlX2ZOyT/baFFGzLSSTRUN5xk4EL0cR/zADnxDuLv5lsY6MU7GegSaj2F2fKz0W74AOr+oACQ
LhK1k3zcOyHAA2V0qe0qGry5yXRSPNOeeoWw1CQOTd3XbUWgtuougfD7TDa3rD/gFxCcX8nETxjV
LUtqo7w1oESUc29n7jGbsrbCH04KWBTI2H4ZRbwpHXc9Xit1ysPl13WofxMadwG0tIrXssAImIHP
koP3ikHVUmR2iBrrkEiaazWKbDioTa3zBKqRla9klExBxs1WoMNuhELh7S8oBOyWY2AQ8K3SMP+H
iM/DUsHALoV8CgwOFJVMEfkojdywXjmYJtcKBHMHnmO1C0MOwhu8HLyd3ep2TJQUNRkWco6QGD5W
2QnHQ1HNl7gEctlJIxOjcasQEJLpY5JbxVBzG0YUKbY0FLjObwRc+oq8BEYYz8I6q88xOBdP8r3H
pqc10yzrVAoVNAYHKGRrE5nUsJAHy++OTxLQPgWQra2mxX3OSE2Uf//ehE9HIP2qqmIsbKm4+oYP
/TtMIRNC4HjDQ04ZZGyQsnZJzJ2nVxUL38JXWg8Hqzb3H3RlnvQ7EKBKJVfqfzrqSxbn4JocQIjV
vr41mM0jehAJF5j7+5KGPw1cRjLNe0h8luW9zp0qOL56jL/qXuZbRFbpBR9uNA0lQUTjjtQd7mTV
Px/Yg7aK9LgtySlqZaciiOG8XkMHB+LzB7fzPE82LOn2AaVjNd5ERVDJrl0XCXkTkDiKa74CGNsq
uB8WUxCkTBOJIRSwfBBZWOt6cEujzb87akZtky9UzEZAJ2RW+x4VNGh9ssJWfMaHX5YJYvkBETWC
IxRhTU0UOHeh1JDpSc01kBfisMaYhIDpcMZQvFTpX0hRRyVtYcI42UG//kptKQAENajGBh2rQ8E2
qWgzx5gRXaZLuO7VMeLAkvRivBQ2KwfZTj6m++9ZIjRdcDEOvtt7Hq/MWeZwGd+LugBcWTyY2tXa
KcTC0Q0BLGeKGtvHp51Zjtk4/37dHpSyFI6J/jkMrLdzSMonmr+a0ETzGXbamSRtmOj8xTQu/KQJ
9A/VPco44W1LiOJ0AIylcOzJfYkM+1rYnrW5GgJe5hSEQDZO0XAd9IMXDzwywcNjT7vukfNbHN3X
tRzBbePNjKbEyXqcLdZSdQ95ecoPrk/xSMep2a6TNUVFKX/hC6pQWVvRGA6JWZ2g0Il9LGXaTHVg
f/yfmoQz0T0qSJjEZldrj1nZcElAwSmEMYmpmzmlRpQtucXz32MGtJSzgcYmpWK8mG1Ouu4KHWma
TwHZ7D1N7blt8PiZmDMlE+x9hW00Hv/hnW9mWIT+kM2znaRPvN0ZnVhFM08yKhC7UpSH+Ww5mnMd
rOh1uF81fvdISrIjifCH2zX/qbuyTi1PfQVmBNe8epP4ZN5AD+GiqwrI58F1LAsW0lFC4SBqAMgF
R76EjpKIWxg89O1e261hWAcrwkrcrg0w/4wQVwlBRNmWJb+mfeZUAKPyD/hJAdpfdlJy8u1YvCws
t3Bm38cy2QkdZe9vVrT5/Jwq1Ibmy8ulQogVZxBtZY50xz/4/LfpEXdCMYWvr2slZKlSljPo1eMv
lu27NrT2I9+5W4lrArkCFXYtETsAH4YOz+k4SLJCxdJ/s4jBVSGfuWMTsG1W0wMlaUIewLWCng4a
cwuUvWMkTxCuOHbg5sc0kRLt6Stjsfzb821WajhcLbAnKf9UgilQQ+YK3RIHwscXbmBWn8J93I2X
Cy9ajKhWM7v5vtJI3JKYWDHUC+b+tf/NkvOyFZOfYluPY9pqW7WU/WmKlLc8iILzRsxnVJSMOiPI
cArWFOWMwDrGubi1vVFpRdTnLJL1VJ8uoJvHG3Xda/kMYjxwL20VOc1XGsKPf9yQHS5ZCTP0L9jt
vgk+biN8E1/e6m3r1vBy1x7m5j4wALJLr6G3QUo1T5DthSD8++kN7hGLbMUuchl9iYHbVDjRe1FV
0cbidwCaVVZvIqE7SW0awr8a0IM7uPdmdMPP+zvRVwYRcR8XJ3oDrq4ysqe1O6wzhxlNWgyYbVN8
SdhDPhNFp7UtTTvmwQwYPM7cxatSWLUJhfu7I5Sa0YiQx687kynvhd0oF/SWkb6jstnLtbzONLbT
HW3GqghlNELLe3HqWPHtYp/p5ChNG2U/dQVAPcHTkBEK8u+QJEqXL/hQn2CK+wAcSGN6am+uK1ql
OakiRj8+t4Qayt3NU+wodD5L9BFOJTzJGwHBDVAog6aMjne/ourmghZ2zR6VwhRQAAqxhHsNfx6l
a3vfI55KygaC4MEDuc6Q2bhZvhlu0tRopAOvO4ALk29TAZk0dt3ckiyBjkMJCioke2Nz6wpik/fi
n1+JXLyw4XYycSY1qcr0wwqA0X0LYGaxOde6p9O3s8vfOOuoD+YliM9wzvy6p5iv1R1lO9F6pZS8
AqRBkxuAYQY+yqyybBc45WVh1Vkku0Z8elkYlcsQ/QDGV2eT5kZ3ZcwBqZ0VRHZklQpuEj0H60gR
1qAsAecs4EnmQLXswE+zzMF5HkX7OMrYPs6+SIoF+lN2aXmz+HQAkyxzMx8/nhs5uYJ06z6auo3c
lb+AutjBjCr8+pKYdN6+ZxeYSrh+sNXg0fAiQto0pJXxMv81ojB19qTORneTGo++0qzO6Oovq30h
HXfCclG3rjbISQ7SMSOC125ihf5wpgUftl6PYDPse84A4VNDxVhKsn6ze0jn+3mutwbUXcsxAOzT
rGOnFKwcpFe6Wj3qI43C2CPHUQCEE3DaUNZFuBG/VChn0eOWQawcygWBhcp3xQ8i3k8LaMcVkYYF
BejKOoSMYuE85Z+CJ36xobEg1edboCxkS1dZGQozptmcClDys5r6mb3FcRIIuthixE9kPlun2XGG
JVZGbCjA85J9dAAKFvdFXs1WD89G2KX0ZcKVTCBPfihNZ5zItvqIUzfv6j8C+IdSoEXx+Z1WAMeP
BbwufmBpVFLhCZttZ0+sorvc3u1SOGfEQ7XOD0fcmqOHHDKMXLZRNdz8mRjbU/oiZRDgO7K4ZCcq
NQ1/8gcup/X3EpDjrTvyS7Ar69vheqS6hNXWjwOXqHsepAQBbUKRtP8PWiR74y/zzLSfSMl8BIdS
0TMuF8pZ+5gflEEqjml8L3iqsju2N0L1VwqkwiCZEEf9yiVbCAspIFY0PQ0V3sxzWSL+ypImxApW
KMtMEkU3lIOyprwi9aCDdmmwnG7wfebVWxAZ5+6KlNvXoL7Ik5IIffjMS2xOnRTp7vtHZNd5baz+
3KPAQK/ctCwaa/wGbwQWf2zFmMGoySsRJcUpNMxrehYnnl7htqSpbyaExuYoyAhI0b2fXFu1Ik+G
4HbeUda7mqnsrlPKkSFDci40BogwSK/IvQF3tqd9YlevNdr1wIIe0j+kwU4A7bUENodT0JfUUh5s
mSL6PTP4kgpg7ebpu63FN93S2iVthlcPDy3UnbHXCPZC8NOrZVgXwwgWOzjUm5R7wBbUTR6/+Aer
R5PmiDbCWdAUTZ5oQsUXSRoedPud14Z3zzBZRpIov/yQrJkYaX3FaagHutQI1VYGdZ21vwQ5+MWh
CnNlrINB9lSAbqNBkBoFHW/QdplNj4WRgqLe280yiyu4880PuK5GPS0rGC5fOFsHb2CSYK03T9M5
NeqGCsiDsf7ZkUUgJm4w+54QYNRcftTeDLMIU8SoMJY+4qShDC2je72soT5amwmzZ/+ilkRJoYnT
RYKRUFKJ2PX8NWFw/AULeBtsrjC+xOsKJD3KLRcjnNR/9J0O+7OfL4mq9AtlDrAy8UaAOvvlXapB
NpV1tglawOXPatgZXqtC8Oc9+czESNQtGQpgyDGAwmWX7yz2+DnCQIoeizGk3MHVwzfR9aZUsavl
mE7CjWB3B7CygPrXmipUcU4PA2II4F/8g0uPsbu0+UfYzh4R1SRWj366b+50cYHRfiIcvbqAkQMP
eHeL/iHLdmINjw2Ou6NSj9GcsTzyfak937hnNG2O+DyfwDNY7Ow6Ar1+qp70IfmSBL34HOfeIqi3
yCp3pn3mSWgQNDBv8J+2W7kyGIKwFCKObZwzq/fcrYQ5x+pvhvTbT8XiXsW+avLknjIEbYM5FL70
VD+LJ5nQ7rZZQlavXwWDEm1Y3kFhXxm1RDpHlMvlgeDaOiP4rXIvUlwCa6di5uQyz/57smalA+R0
YN8fMgSmfoMvRfPdJNPk0PX0EoaaUV/LgcD+jGJG71FlZNezemoTS/sls2dJROIhSbimXkwWp+aE
SZW6ycJpG+6VApbWObJWMGsZB8VIOUHG8jatOWMVwdN21hV7wOd/537i7ttbFOV11imbd8ABqLuq
If4l+X4pwEoTMI7qMD67ilc7a5PmP2BKKYK7i/Ng4FZNA3H59jYolr5hCIK/zoXwlQtqH6Tg3Iee
ckEcxdrKUAzDmmE9gv1gEe1nIstH/EETUO4J8rD9QJw55ko3688rXBnZ8IGzunV7xsYKCkSmBtzX
8yvQA77UwvtrH/4s0YRZwhVf1m/b6W9mUSHO6GFHxQFT+dwiHv3zwdb2dRUzCG4bmBCEJKleBNuY
wlr32rGyuKSwG31E9kn63VdlCNEuaywQ1Ugnxg8rnCCmq5QWlbViMoxfEZfE3BAJdpuCix2XWQJD
KZXBQR20REAWsbZ1jwc0xVjbMnife3hpX4lx/kGSdM17YbvkAZ4hJwWuwnIAsmMBl/7AZ47S+8I7
2FlIsJJGkbJKuiiDPB1hXfSO5z4IPLyYuYikcCdP8O6fjnMuZjAeT2wGBspxnaweKrW9PMJ5/wco
MiZCyGY7o5myheVuPpma98s+lpSnQinLaKXF18ZOwTSzqKTrdkaeLtmvl6dp7jI0SbZzV9RUt9yD
3LLhCvo6gc5eeLaul7Q2iIO0FabHOhZg2ytGalytmIRHX0eicZlcf6z8OEJeucICmY5sTcHhaSCT
eM47SFVPfTzk/0rLxZ5v25dXs43MS5Q4rqsxj3PWzuYd+DeR61AD9O01Yt/HNyGCiiPQQeAS0VxR
LeKg7xUGBblALF8ZT524754YquH+PnM121KIBymMQEc+jpgLUHwC/OtzCbRvh0Sndv6hwq62jX/s
5+3KDMnY2uH1OCa44BcqBpigmxpLZ9u1Z1j4iQWKHE1putiBQxaVvDFzfJi98lP8RfBWDqVp2uvC
9knb0oHZ9QZd7UPTNP0hKhSMSjvd3EyaPVwPYAXVsf4ZY4jh1U46G1WKmG7bj6lH8H6kQyxb74rk
iX9dQxlBJRtfkJIq0/PMHZ/rF2NuhJueMMOzvl8Yurqe7AEjlIMNsF0DsHOwiVj5OlsUPi70TceP
JJ8Vu+EUj+CVtqzl9WDeeV3ZQilA78jys/zLAHXmIGyONs6hVh9wI0+rFv2cMV+IoO20U+9D3tbg
I2ocQw/6VejeT8UEl6OlToM7/ZJGFuXTEdjyYysm3Akpe+WXqx0tMPw+8aV2+UhoNpV0B9oUZFwg
jVUlujfTnf4y0VajHsZaJGNH983qHECeFHzUOIP+0h5e1fuhJEs+nvGAMCwk2dn56kZj9MLNDWYs
Qxwszm5+wmJ8F2AJTb2C+f8w8c/+o23ydBRaN/d3+cMZtfVcyeycTaROENewwfLI7Acb/G3LJYdz
gjthWlp0gyw3YaGQsFQQRNL202uv2pPIPTYHvNWEzkVu4tJn2qmVdviSkLqGlIGdv8+E05H5Qt4n
iUtQdy2WI2GZQAg/dTaSyKlwKihrO3YvrdbYA+C/atWXPE7BtZCXGlvSJ4iBVt4yzfzIZ439zKT0
nk+XvMMei7s/jsPrqGK9hSQSd3KiC28ES5BrM1ryUqvpoVsVTALbkxYD0La5O2RwapjQ2aifQm7o
6E9IjTd8dkIxLm5sWXdda5++G1mNIAWIUiT1kX7JPB3bydjCBVQmuokBPAIUGEFVm7YbYWpZe9u1
j1WOoF1w5uLBw8RVSGTLUNjamaP8P55FkJaF6/3ci5AHvFYmnMT95iTyiUcgNR9F402NHab7G2Ve
BfWiCaH9b62DMAPN5+3D9nNHPgdJeH+xtUp7cecsqsbD2lyZZSoDG0KybHj0dSunglgmY1l4Pizd
Y7OKq/PaZpmKef5YwWE/PXC7zPGLwKpR7HBsaPauXPDJxsE0S8VV/LOlJAFBpAEFxZZMyQQek0ac
xgy95NPq5oyme7N4fgjRLQD5PRw5a55OVY/FVF/9bHnMc3s6Ls0/uj3H82udbJbwF+lC28BQtR7O
mzzTsTUmqtSZJ4CeOcSjNmdq5Bq1gzM3ARwbM8XoK9/4OTxN99Ach1nKNYfCNRkUEuooet2K9/dg
HfzTfr4psRYWtW4GFUAJpIZMam4ZgRAZCCT28ZVCumZjxnH5v7iCsAO/e0dWDytbPTT1gVTc4430
zuwITOunfyW9eAjGMijqUUn0G97R2/9KS/UqPc+CTxha99eA0xOgG8cy1Ok8p7fakX48pXGrTr2O
cTVa+EDBFSce3nBNZhPYLbPj/y4w4aJHI9BpctStPp4i1YAgWW+e3cMJzTzo1cpD96TlfcLCWAmO
5JRjSwQSPkV6ezGC4xIgzJdX5LzD8fTJR1RpN3alHHH6czigCHsz+9rMEKOKTNyF1WoM0q3G1qk1
QUeqVuJRYukbsQARvYOcTul1LCfVh0a97j1xrmSUGrF3n1MBLrDf4NZTttlo9ptt8ewqZgLBg57m
OBLDEBaveFZyAqdIpWWBu8+r4iej07E5psx4gto3h5MwrgW5NuuU/PXRodrV2WlBSvIdsZfQ+Jzu
QvZbMiCxbZm5h2vM5buj5P5kbJ+jTvhmBxOYzXeC8MHa2EZQTsQtw/zFAP8z3vz3eSOqOetGF8Vl
5hXg7yruwrsdd9Ko3tc7xuVTkMLHySE3YFUShO9yrthlq0wBmJKamTAaja7iiMBHdrIMGPm9D+p6
s1VA9pewhRbweB7zUmStn6RArh7p+DD9pMOnSsaqfsReujXgS31js3JoB1wEClq0Kd+ybH7BiBq0
Q3XERhJOI9hU7bblFxzHQYr64bW1RYSj9oW2LCtMvlfr2ZBdf3uBMxFULltNa5igjQhUmfJL3OAc
VwgJPx48lmJWSK9/pZXsKhuhodKR+63i8fFdJTQPDj0DO36v4LVYkpAf+R6I4DbkHJQ7MUuv5bMN
USAAsst07qRUmNGcaN1tMgJPN0OqBufD+RtsEO3SvzJFh4Ytk37d2Jh+FkG6KmOeihgB/iWkt69B
nrrrID40bwip5MvygL4iGQg4K6Lk1YjtLg/0ppDkkhOUayarGhsLVCTGkVIqwS/YGs3QI5WKmqLK
081NqfgpFnHVAAe75M37LDfT3311Yl9CsRu3+pZUxyDaqgqR6TVM43Qc2ddR2hyWJP09L1VU6K9O
EtEt8JF6A9SB7zsXHLQHRiaRgqyKZJRpz1lnVywQ5uKhv4RMMi1mps7BCWhurUYT+NaOwlMLcdal
VZGxM2Mp2B8oKbiuOFWmsKNkxPeym3mS4u6oWaFBSsb3pv/DlM9ErcNWIO55X422QYxpRfcQSdHB
Jxqx5Pg2EWr1oYHUIYLOPfr7gkq/vbJXs3wWAmkilznqm4jx/3x+PxRuLKy8VvXY00P4P2pvzMgW
xcHxXtJS1jd6zG7GzdVOEKsFgmFQNn8P9IQRdrD3B6mZM/XNjcZZFEezGZPTw0X5BQ+iKTWTJlLw
tKspyU8acuWDqEa25l1NZWCATcGf3CF+FKbEgvzAW/mDING+b9ut0gzEA6k87fx6mXrheLKZJL7v
H92vmSEBa2w8z9keY3wCdWoTyynXqO4Bhe64J20sjqd17A/aet0/MjysNi+Fwu3vdFa0VTwrVlt9
c71YYt1hz+jG/z5C+QjWwitvvR47Ve3flC+6i6TkneDIIitpEZAAteoWpylqFUb3E0jyR3t3mAGX
mBfv/NZIY9+C40EK4vUoF8B4iWxPHVO05vzAgrV1eoDhfB/GbiL3FAHK8IqSq9ab/FLq98nuDZpY
q/btrW2J69UD5Y9HhrqpCtse50l7xoi7XvKKbQkqTkuVFx4uHis75n1A2UvHRYjVbMePPG0++CKk
O073Y3nxB9c9rI1rKiOPJbKAwGnAoYgQvIo62IzMiaE9vGIQT2iYVTrU3FFQM8BAAqTZl79BovLE
7GF2WENvvpxjnphgQhSGnzHgkGq5EG9ucV20TPFhyu23tPdLg/5FJn8+Z/OviO/CO+xEz4yt6CkV
XCM4e2WdWQspWzyhTKmp0gjMMMJA+04hx716posbri8NSkWcqaSxdfZZI5pdp5vIUzFiNCLEdGDy
xqzToVCzvey3GNZYNmTrym+BkPm2AT7Eo8plhAAXNhw9QnnrA+V5L8QZkoB6qmi8T/vsoIcrrnHy
einVMaBWGQlkodczBlCLrsNdRnRKyUNXaDZrxhEx6IkRuzN3h7SvNqWuw4dynSBnKg0FcesaA6D2
bvAu4rFWd578U9ZSdwu0GyDjBhDopaJW/4SJhLyOydh3oNc9ecBVDnC69utCumm4JOyDw2f3lljz
OwDS4iNNMY7VWdVP1wAFnULl1Pcm3Jc1goM2Fa9YylLzGUbX+bCHRXdLtQ0lQtOPCHEg7I3kDPi7
DYjQ2pRF2yq5vZ4HqCs3HOXkU75CqkgnwHqU1zffYK0E3ibuBovM5KgpSEwNYAsKyvdfWqz9QJaA
EoSkxPYSTyyBoa9zxqntb4IivI/OHvix8cbypzpe7dC7aUH6ZowJRryvlmOCm6BlLOoGaya7g/Mb
CDs/CRyWbdYEAxvu66hrPF4w1rfIJj3RxwIVSGmjn6QfCrHY932uLp4HtndfEm/Cm59PDI+DEiAa
fKqqin89/N3o+BSE+K+7GXQqGS9UnRHr0v+07RpSB8LiXHduKmnURYMh2pHoXIYGWd8GEUErJAm7
cuR/GIdOfWhuYg0t0FNLALmlLwy8tJYCkkQcPn2OQlsWobPh6D/uhd+CB5Ex0bFwaq/YKJt9osbU
OJ+jywGG0Y3y8g4Y0JK2xJecohTdNyxeumsXQMT7QqfFJCxKcPZ3oX1FyygxxIiGqaM3iTj/Gywb
oSKvshtoN8lHCgkN+Zn9n1kU90Vln9a9OF7qly94cRmz8fQaZg3LWQ3G2j31i6j+r3uy6h1VWhnD
3MOKIEv1pi4BqTKLFx0SoCEqUuQstAYVUlESfo0VoC4gQPXQPDS4lv1Mp393wIVi1oLVRR3yv2WG
cCDoEIhus9fajewsqLNg2r8lI1FDrKFoNjHSpISuLzpiJt6k0XAH2i2Iyio8+0MG0Sdluvu6QmCT
xfY4CmKJlClcmPV7OJ8D6KUspCNEVfh6msusNeK7mxH6QXmai+uKXYPovyxr7iYq5aK5n7XxBpjH
NiihjLc2B/CiyaPBwXmVgLMAwLskeveo8WAQI7P/IsZ8sPlj6inZh8G75nD8SUTd8YqWfuiik2PE
0Lc4YKB+Dw20VTy/umfQvMXdmvbajB0euxLlgQW/2ds4v+zAoMF2AjjQ8CcPQQr6g+RyIaCFbvGF
9UezJ93e2O89MLbvyDVd/ICnx9/1lMJm6+QV+DYqTqcdZu8Sbl+NAi6K2ucn6/10QBYaN8tfVM/G
nMIg3v32Q4YWSBSsgBwCYQ856yk3JlJZQvRSzWkdDBZqerPJlujYAUHF7izCkV0QVQXHNiJzPW0z
85BdRT3sRvvDQiwMn95eJTnQ+gWtGJ6s6Gom+Ug4zcNd8zupTVpaBnicS9ovEqtdAWhr2VQ812A/
szdfdue8tic8YRltu+cNIS/8JfnxK7cwqdUME6lrtVeFPM/Q7g5Y3W23iE4mBjsNskv77gqMKESH
M7S5NSvlgqV1wHErN1051jgHXz0fpV1GK4EUEQWvQcNwACWBGsNOdRrb5hXDDZZRVJzwfpnRI9/r
ySOrFNGLv3Ys0T+L5JtXhrFmlnXQ79G120E20EXA49OfCHRe1EjjmiKRp6mMub0+rGTQVBVcSHix
tyx3GDILSAiGU/x9/4DpIIIkMIvzFNfmYprlXTqvYRSsM8APvXhs5OjP2bRK3AzCyw8bz8xF1Z1n
9RsR7sPoMRiUuFix79hMt8zYakAwaj3AgoJxQULLvBbitF/3VpAJJV30iFk90pXYWcjbLtGp9SGc
brUpQS5R0JxxhuhktzetHIWlI776J8eD3lTp758Y30objR2THg822fM5Ko1ia+zVVPNDgPGIdyVi
ssGINimP6OlwYMiz19PtOXFtQyQ/KnoT/cNxgF9AcfJMA1zZfCk03w/dPUQtzjOPwoaJKWTgyEXC
3EFOLm93u4uTOE/EYLUHNm5A6MRGUxxWtOk2BTCBE2HtR3m0Z82L6kdJ+dVk4YcE9lU0r/4i1k2P
V6d28j0h9HwVrpIVxU+xa57RznLHuu/qCyazocrNCQLi/CTk/NmdGdXG6kDMKsQWjm2fijs6ZbQ0
v1HQmpVOAEfQQIC5J4+lmHEHqtfM8Pc71naWFsN18POJZvuyW06zughbqtm/uH5ERXSahCUscXku
wAA2tsUm5QtTdVNE2OTVpZ2LWS0jZs079NazABeTptExUahZuPICj4Dh3rs1CsJ5XmV+HVFXV4GR
lKSr/WdJGxgE2EO2pF6vF70xVMheQUiRd4WjLxnFDSYjFa8E0HBOm01ix0vOu7puX3WXNcKIHKhe
lLRPaqfKQ26tPQQSiDNuN3oRvgBZluK1mNfNlwl5Ku8aMbDteJmklGkpLQGH+VKN04p7xCfwsKWJ
yL7juWn6j5jmaUUNFt6TT5w6suXNDJEYlZ3+ENg7ciG2HRonvEoO45OJuPUCgnOMTH1c1LIi6fa/
7akrU21doBXOKef5zEzWtEf/zvJuv0G8mpAHhVelRlAEAH7fj6BQoBWcFgjY6TewNnf0fx/kk2Sn
XtSyhOcU9NYYd9qSQEMpCRTmLimp6r2u6hQ8kx8edtsIwCK2jHuaEvSUQRB3a3nkCDnWzAAF9Usy
GQfZxAQfqtLPcjIT93q9M8iseh/AFOqH/z4HppzxTvKCrOqW9F1MKgmXX279sMj74uTsAyZmvNWu
aWCLtVqEyjG9ykKHNtOysjNAhMLqBK4XPC+Rl1Ehg+6AqhoVoGR6Q9xvIy4XZWJzI2b/apEADnrY
JmsFLAMlrPghYFoUa6UdHL92GZ7ZfO7vvckoYqiw1fhHEE8gxTVY1jMR/EF+2cQCfTbJTWWt9mEe
4i+h6fMddm6typNt3eer2/j9kmkBwVWbVOw4ECLEtS8sqCJx01hsIfrLMk2jxHIdfmLaeT7GHEip
1KY7ttPX+BV4eiXIoSS6g6EynEVRvXZ+L+GR8ZjxMy/cbegayRdC5EwBrxJ3/pyxbPUY8EeF06nc
NqHlB54KNfNI+rlrbiBTVAv15VLST+y7rXcOmHWHXApzk0jc1K+/3UiLwvSALTXgrRINpSRF9UMH
5TjX460nz9TZQrsdh09b8xnEZpoXWqDW3OLRONfoP7GIWuKHA+Km2eWXDBlGJoHcJuX7fnqj4h2g
uF5AkKk43zyiD+TnY/+Rb0O7hOVm+20FUTCiWxnZ/z2D8YWscnG9mIrO9jh0qYHEmYU4c5N+c4YY
BwQmDOvG3/D48hNmVXMHB35UgsWk1l2INnL0jPCU+pqjle+qRuPjOeqjifKK+STRDh1XMc6ZNA0y
olnczDeNsHHSeMKA/xtthrV3ZePrDyi1JxLokpRiJRhfC9kNHxzqAC49jHUxZ4h/U5VMqnVXXSiU
h35F0lABTnQEGs+Wt+Y7awyLcYi++3Yz8rbHAaU1OPhn/7RXsoI/nKCRYR9i0XphBOiMUMb8oaWx
+JxL6CatPR0X+cAyA3RhyTpXwo9+Ym6k85b67xVez+wqKO38w0VWSixHygHGIvqRWuzUofsYh1Nv
TkXrKVH38EMmFYb4HHKdcTmOHTCw5GEIDo7+kyt8ebUuQKVclxMsPVpfUgpgKZu0EDEOmazJuCNv
FWZ9BP7e6ImV8G1hsZ7vjR+H/2MyV8/X/HWbfrVfzSaC8gDtjVv01zfGrqiV1aSVgoWuqm9XgJht
U1CqDwowmvIQHraCALLCFuT403zJ+pfbe4Y4C8peQgWH63+hm0h/hGErj2uHQtaLyNCV5+KE1z9/
gTxLozeZtXdURTYyDuhJwW403mXrzoSWBKZmptA1PRyOhKQmPcFzYNM+0VHSsXf9FTb/3h+qUT3w
qf/NNAmFq0TXAK1+DHjuyuBILqO0dBlbAOzgZ4/85lYzTF4vhlTeLkLKd8GdZiYkHudihBtYPNuv
lpLpmxVYVJQNeuNjoKKopCnlbX1LyJr7bF+MvEC/+V4b67cuMxcgqNadN4Xi7mPc0Y/vd+hpfp1a
GYeDMU7dx9UTWWIXH0XIIqfYP8Ce0EabFcojpX0dKZm1ns8h+NfUZj2RaCRVyK028SbvfwIox0jl
ErA/U/enO9sjyZUaRWhI4CB5FuSMEvJ0oU+hTetIGqSsujZfZhhFGNZO7yq7s2HW40QIKOv5/9ul
mk+imcKbL0NUL4NBZWfuSwkLb8Qp221wsJn7VcuxQNZ6WT8+rpcd5XB7QR1gwmtbI+Bl6ccUBnyD
o6crGUIEt8i5c5av0DRjAciFHgXTOGCjjNIl7BTizFxxAohduLUyyYNC0Iw+odwFOMOCn09spHF0
mtDCrisTrhapzvNIb4hbXS6aDs7rTEu2Hq3HyfpTN9Dy2nZ0hVrBZdqRdxXXSpCOTIScNkN+4pmZ
wrTACiJ/M8NONV6/54QuLutyWu2+XQOybqGzK18Lc0gBAM0JVRZGxxO0nb3nFagkmnsE4nuJwSur
7638eIsSbr4qM5L3pU6dPkw2EM+hA+zIzYvIFZ3GHMO7AiZ3IEfv/SUw6jBkkxvoZAst283yTq/9
wTG1UbgxKDLtzyyOzO0cJJqbaIihtKrrirVWi4zYHxzLIl1ZKjs491uw0TtSM/qju1Cz1aPAMV5u
F/cxO+xMxalCXLBlaxHkKQnOAGesTw0JO8dq0RykKPIcR5SN6fOtjrNySrHl90fPOTL1jVbmHClu
ZFznrQ2l/n/1aLN6KyeG3xX7/HA9y7RkDd5m7+Z0/lopQcVjn29jViy7hECatzniPrOYoCH/xPqL
/UrcwoJ+VfXMck8mnqYBjWO7Ib+EAhF09ZlWvNl8OfI4aQfSPd6aZQEpM2cRLfz8tPsJHBNLOsy+
NdP5ExNeeREcrlv/pf4aY9EhhrQCsTS0+pLk6kClaPZpWfsDRAaEOrIfGQDzAIZMaB5qMa/9GkaF
uKm96e8spSGetfbhY4ON0yDhFN521Y7Jnul7geiv0Cr5iH2X0DEhSVrIddSuJl3wpHLhv47t16aT
uLCXdU7/5vKq8rzj1Bn4wAVGryvYYer7r3ekuBLuO+V8eAoFADBox+kB6vwqppyPXgv2078t5cCf
6AVD3E31UqDbnyiRKLwahvHiBLzGztnGA/V16CoYyecWVpik8qpOh1ppzmym5lMRv19NcR1/BN2X
p9ydzd5soKvpvNntOL5m049Kof6xgERZTreItMHQCB+LMZLYOynTJvluyX6bKM16yExvsCk6yppE
TVsHSRZ/uoiWK7QkCzGtAefytX7L/VagRhks1e7VZ/rbhesjr/BLWpBYAfE6OX3xXkH4spqG3rmd
hUuDotQ6WDO7yx73DD5yPmytLhz0mENmonIW4QnLTdhA95stQLin5/dujgpIINAJJal9p43Y42WH
uvYdB+D18uKXC4E0UCuF5XhjXj2jG91RyUZLcM8Vxgq2ssOywA+lXN8ctC6CoFil6gbTJrJ8wGV3
sxPmaCsuwdZCDbJbMEnmEQ+GSa8mdL5Sy9sh8+37v60X6oWp4f7GVN6QlEuxlaV65+x99XV5Qdcd
3gy/zUBtZZu7hUJdnu20lMOzYEc1idjc0OTQTamom5+3jjp+XUF+6XqLddy1b/ES9jVBLZITltHz
JTTCrdtJkO3GDhQyCjOLssW6JuAJZGzsi5sGx5kDTRmi7n+mtCjF3blKJ+QbkmEqkN3bkUfqp2fD
IpEOuNy9aYRz1lImasvG8J+cETsRmbJRaT87yZbuzpwRLNFqinmPR6VSosJDQ1MkluedPoXjvFxl
QLM9zuyNgPAYjEiO10ltsSAo2NhvT+VikYTTvEpaHclacsMjk2lI/PlaB4iwpiUw7jBMQeDAh6si
RE1fieo1N2ox13Wb6Ls27unwH3GShzKppbr4wXtSyJ++FSOwFzy+vGjJ5kF3G2PRapZc49fp0ZXz
q3jkr2T7GYhJuX9OjNGJPL9vUIgP8+DkNq+C2XZA+Y1MIwTmyLgp/gbWVOp6rn+fklpFLVfmW9tv
lWlfZnGSolRwwPSN7CDly0gooksaOFCsTrKvR3MA3JDIy1HV2+R9NAR+rvoLYM1y0I+NT95bUXh4
yRAMOlM31bTGjnRwldX2S7Q1t0Ekkop2hQ8twCpdcsDMkeEn1yjd8kcQyGvh3H05kkay+3IEA01o
PpXUAADmsolG7Vqo7TSALhyvnsRwSn90vz8dS5qYNoLuCYk0j8rUbYFG+KLUDjFY1HXQKfsU7MPi
uhY/drR5p/8n6jbBsNcf4YCG0TOYi+bICOAJrJ/wCKSVVtfnPbYSF8RxEWGrdM2Td/By072YAd9w
gBXwuPw+0ybme4ZYTktuTGTGn04yK248tLGjxnsHFZxUuHdOFUY56IX3R1XWJF4BllrhyQ5DMd7V
1I8wxVQa7yalXvnTPjDEGz/9TyrbEQpBdHnCm3zpNIBwcBww/81v1UJaMn9PvJSnkWX9ghiQdDRT
pQq2bmPeJLgwvrQbUCNQb3BXOYdWuKaTOYoWTx25cr4yNzI5CbY0CnoJYv9GDbQhUaOWNDLEW/O6
TsVeKujDknisOVdyQRynz5zG3QcUAakLENmcOUcVW81dyWjEdL967R0NXBwbZbUQOKwalOtuHNYN
G0UqzVfNUI9ZyZ7zW0K0KTsNvA1Zyzf0qd8mSKg/QDLo55E34bLLyVs8+//g0RymEzJegLxM6Hwy
WCIy+UGaP1Pf7MlOoPA4AZpRYvlZDdg+Nnp+64AxGqajmKs3XorYEW59zEhf1246z1cUahR6O1JE
ZjhAnP7NigiPxc5FtAYupk+OMKfe3MRaNmouHUi76i7qAJQVj5oYX9ic2YHG/aljaxEHdt7QaiMO
zH8atmpleE8y+J/Ul8eZL6kDeOnTEmIrlptFTLqRT3xrmIUZR/45+8wpxA1/RXC1HSykCYPprzfW
ejNf7sF3UmtVdIrVWFFEyu9T0GAb8auPm/05sMB9dVBr+7yBVXB04q+q+HOGd9LmAXo2s74aEjf5
ksdSAXKZoNwvROzPVNhu2XBrGsjbAc/J6gDZqDy8QuPHmaJf5GEQmxikzrUukawpw9DQawzs7prG
FBr/pC/YZJdssUvCxULtMbQ5u4x3CEnmsdVjU9Lc1c9O7EGIvzZiD9zGzkqw8r1cnUS7OEjhV4V+
SmPDtULdJHi0X8F6TIBkLjtLcFRyImj47T5V1KO66uHJJCwILcGuN7A6qlV7PdxyrIloBKFSJhfC
gow9JyMFTxlGbAUag2iNkNN41pebhXin/Cvk//aewwgXhs9HmOsfCmRAb+k+mmce8SOFJh4YEFfe
npDR4+q1jKpgFNDxuj1ovKs/xSIfZj2ZIjRbeXFvA8JBpbR2c0GYtqTqkigIraAD5xo+6tVnBwBH
viLxg9QPnUp7WYkfIBCxD4vVmRxr+/si5P65JiUkIZhiCuexyGd+jVRn1hE0aHk5x7v1n7gi1rrd
JAmJSc1jkj9y2LCaE0zTtnFgmJZ02t4ZN/gZwW2Kc9SNVlfVyb1eddDJ92ZW8nxOUifYGgsqinoX
Q9TbiTxncSaOAbvK9hIAQzArZYEUFsW/dyz/feSsZatF3eOmlAfXaP1SZtPFM0E3S4MGFeUwbQlB
jd6ufjLKZ21FK/PDNPelmA0tb2ICJKxROEmjjoS1wZs5Tp2x4EG+92WXHVuk/h/J3nig8Td7Kmwq
pugtiex5/nBRFncfsMXMs3nDMWtZc02387il8mxzbs58bLoi1GtPi1DBQWGxW2dinFwoy5V4j5Zq
N+mmuGzfzHE+/sgI2zGjuBDOLm/OokRLrYpx3WRBNDfrBT5R1sJRdKBs6De5LXd6JEZ+9XK3u2UL
c5Z4Tav119uz3cNX/nkiZ7pEihhpjQ9IW1M74fgwGG4wb3tqpzekG1B5rCL5p225CDTC70cJgl4D
55/mpW+WVeYI56PwYOjQnzMv5bFQuewr0xkA1l6UNlIkDcj3PxTauVSS9ioGnStO41pYOnEcM5ll
SEuMldjEqKtgFSlDljnH38DUQWU1S92UKyRI7Ng9Cu3TnEN+cRWwLYsuiyy8+7vJqheASBikqmn4
FhChM2MpNPX/zC/XHjZS8xqZ0sQFUoPG8oFWRjogWMIcN41UhC4A5bQpUrh7UGK1vI1r8ErZlphq
JOJh4mTK6swCkHi7jVaLAxEXXeGOcx8vgM10XEbZ1QGjIeLVd4DJZqchMPdHcqYx87cd/6Xe3s5W
uiLGoFUZOoXJGj3ADiiYe83hG+2EKO5malGKKTsITOUy69CR0DO+R9osPQwrXkGCS1UPtAhW28mZ
WlvRH3+m/jdU9XdWxJd67UCPT5Z3XZnrKa3dBR0XqH3O4vhZEDKuEe8IjbiyMdoKIpqo1yN/qztb
8IFCdy/7Iu0T9rAb1G8DZ4h5myiOpn7yoYap+fBqZe3zy4iImUu5TBaUAIh33xf93OzuvxAvPIkf
C/qSAMcEHiO2iHDfpIfPuycaH5wV6+7GVKf+YsNFyfaPyvx++soTzz1TEkPwjppJGie1wGTMol3u
HX8wnM4lVtuNDb0bLXjdYkxhzSSWCc+JiGU14Bk5ypRJ4acnXkh9pPRiLpyGvfDqcne0kIyg2mfF
m2bRRPcM9VFjU2+zB1dy9zXjJNNzCxbrf6pf+iiP8Y3mrhVBL00CsVXWfcHOBvVo6zdg6MJKUhkV
H8mCiG5VH+qGuTwZzCFKTaUtltq59xoaxqLlGng4DbEzR8WGJ5mSyodf77xtEwPsjhCdV6C4vxLb
Yz3/nV/d+6ls6FgNkoJXq67LMrLzI5msMGhcFyBWtGv18INS4BVZ9aV/oLuwPEFzC+HBBDL8S6VQ
MpqRGvj+hK2kmsM+PNG9/ZfbJ/V7vXUEqkUjsWIctTmF/NoHUzYai9tVTA4T3vlBQzO0B9c3SIri
zILw28nlT1jea9eQg2t7pWMpdxoUkhNeJNvCxc3f7ob2gP2RBhNCOuj97Ls6vJj6ZdAkOs+v2tRg
3n/E4leWNdQX8UThj/7X2BRqqoDMQgzL5/m85eJYKCftT331o4wqg5SY5FBZHjqAPxkZIZKAD56t
JOF23G0z9ztQ1avWp/m3m05MUC9hzpxYewhq+16CCN3/IfHLRWXiUiLDnhz6pk1bmzXCONGMSLoG
fn39isA0q+zFmQBVRtwSdfhmPJrSVCTneRxPZ+mbqBnkvZbQ9rXcPO3YBE3bk7YWvSWV7+jptm8B
uaU0bxdRJE2neS9cpu1D2RYuD9Xw89On5H2AGRB2ncl30hhFDr0fpSmAtA66x18NBRmO7PMJL4Cq
+pSOXcQlTEeT/BMiOGZLDv+tXdThBgUevSFQL357723anxwK+1y9fARLXdMjJ2zkujGpYomP1/f9
WM0sPvX7rEAhNbenyfQnu21eLnT3vwrrh8bDg77iKbj6Kp9XLXS6g+rEO6Itw3oqOyuPCjL7ouoN
0hzEVvDApMTsz7fFxmVkIETMSs/O3OCqJfR9Yt6GH0cLtWLYb4essJ/uECcy1ODEQYKYKGeva+6i
IkAyd9u7O/pHM/jB2FMbnW70BInZc25FZ8I//ISluwL7w31vLlfqyPX8RHXWu7eJ0onvXX/IX+79
ICJW1A8oc2FFiD+7JXqyEOT00njozb7vSpAEZTeM3D6TPFMoDLA3o/PAW1hlN6ZmrxCBwcHECqRn
tfC/18p7mLcmOQeoJ/aaXPPnsZVi9l7EvbL8bX+nuBCQbDP9t05U8p7kf/P8FblkYDLN05PqkR6O
g5um4Oxzjeh3kCdZps26Xk3uIO9sYlxFsdse10oMzASSvll/+ttxSW5yZofxL8RozlCdec67ulZY
SdJBpnHv5pLPKk2Khg1Z1ERlojdXJSty32gAV37PEyZ9QniPRBkdfSkTkmBKdLpkiaFdkxopwXw5
GjjlzU+jnhX+/5vDcM6DH++E0/YLWLqTaRpUnD+Ukdd2BVtd1MuCxUDMVtZ/z45JJhrNmZEkq+gx
19hw5JFTMTRztCRQUzPQR/fm1oZ+mU/SKgjg39+gXsZt7iY0hns9wNiHiyedUsxABDXpZVQ3upTp
xWP1rAaQUnZo8dew/I8sYiaC6y3fpsQ1iLEQ8ONM8A/1XzTlIOc97rC5Z23e8YfSshZKcihHCHlD
eudCx1OigRhM3+5ZJp7++FuE5A+z5fROyMKHgoKdJ+zM2n5AprH8agmviQxSvl2zYSrIJwAeP9KR
ov9PdmVTTChd1zYjek4Jl9ytqiVgfThHCBOgk0Gmfoj5BGftBQvNFSC6xSq2mFpBVncNZD962pGb
3/iUh7idZMKbb+msSP+q3B8b/qvKcDMdJTLVAU6Oc4QHNZxP3lLv/VUeqkgT8VXI1dhQHRjggLmA
jl1MePbXV9+5uCZ9ffYZb54ZAPeVi7fooa0xJWq1TQFnZzzA41XDVx/Psa7BjkvmADYGH59mQpqb
N/nFu0jdBZj6tHha8+9LYH0aAs6TbwHX8KxxQ+QrBSn7oeXFt7awRIiSOve2+TAnWgB/LEpL4IBA
o7406BK7ZYTW9YKKmSQhuueCkcswHmugny8Z4S30brY4A6p1UFjthK/H/1/edtY1myeJPHqG9gmC
xZc6x5f0nVudB/Tnb5ut93Nf2W8o7W2rXjXYtenZ8oumyib0aAGxTUf9uBqTg4CRkvjGJtyvF39Q
+C8sthma/tc/r86/Bcctq0Wa+3HynNDPiquGJqmFrII+cwDIB5lP+vGEa1jUF3kS86N1wt1jS0XC
TQ/rXN5B4spkD6gKkJFevwnxaETOrRb31V14Ywut1b2KChuy/GZ7TEvTrg6qg60+xukYwEy49JZe
ux8YAhpUCdIAi9AaBShtktO4eAX8ZE3fFBThZQyTn+ihNHY01+HtcKEW0omU7oSgcx1uL+DicHBe
3K0mVi4bRqzC8hHkLriE45xGpKktWG4hXpoAhe6X+/QAEjAmcqdWamJ4iCMrQ8oug4ImK9rLgvVy
1wGlAptdunaL8HHKytJo/B1tueuIATxqgLii23gEhk+dhBtjTJeLwZ/t24R7yA5bWe/HRPaZF4jo
0L2LKHT7bKRgT0Mennc95aOCkrL+kLMGeNkbCK4ojd0vDj2rfZZnYyfbdaYvF05BhwqlcSNRY0cS
WfQKEkzhlPtEe/Yal2PmQI5ea9t+w2j+tF8n44OfTKXMRdR+PV+8LJbnIOpYcryGl1VqOZ4y0i74
3exjJiv5MpCKmGb/1VyHq+hATqpL8fEeQzhsbbsOKKhJMpChLwkuTsL/Eswul8v4LsVJZ3mQqMn9
hWyhbAc9cU38akjAIDfp9jsHYu0WUzA2fewmfA56rlhftWfcz67WEkPsZaWQWUr2CUAMFpQCtAB3
Aw6Ma0Uia+XcYS473Zz7HS7AoNGmVh+9aeqUn4yGQqPJ/iihFLDp8IIJjtdcbXlk3AMsDCNR8Mye
RK+wIMOyWk3FBJ+Z0+T553T3v8Jk0xi1smZrDN4l0BcLpd9pGdxJNziBoW9LwqHogJ6RtPfdnw22
Zm5f3wHuK/k6VAXR141HN3y2RG2BPPLDGH1liZ0cyAdNzM4B7KU5UnruBs2nkOtBeQBjRivyhJ9N
GZk2HmmoGiqn2KKSARUsGI45+0PuuKReBpS4rectly13qIQtLPaT2RIY+/dhhgR+g4PU2NS/mQOQ
qFh/CpcKYb6GApPSEThlt4NtLFdiFDnoLs7UywZ7izFeowvNzXk7OHol3RmYYFcZwo2AhIIvUfjV
MOFy8Q2SdVfWrskgzUpjrZkdjWK8Fqda9EFpHE+xLvpV1PoDArMKTvoO/WIXAH6EnxRb/klAWmi8
8HKWZeHiXRZT3M+jcWDxh4FIeNcp2OHgxhdTGG3vwZ/DXe7nBvIQaOv+99j8Os+EM2T8ld5j7Zyb
SlSg4awNRKSS4LVylUDPOi5Hp5csB3fgb4M8QdEPzp9sa2YWcmRBtL+0Wg7/pmo4rGdptTWL4wfU
OhHgPGAErWO88vdCPuCc1WZnYCk9sECyIgzcxRTW//1c+scTd1XeHF8cP1vnrY5KC63Ayr6EKiRA
FntYW1yv5x4W/hw0qKD6MiBkWXjzPM2Lp7AH7cuoS8etbJ77qPFeZisl8RVh6j7FEe6Q75xX29Bf
0VFe+4sa4SUUh+DvaqD6iX5s55qFESFAHKgnbkj0jEZilbXUKnLjecN3xavloqDEgnMU/sdK1f/X
s1m56dCqh4bp5tpv9UY87i+ahtQa+CrUSvF3SiWDlOkkXdLprDGGmNUAhn6jyoOWi8gP9Rb8vIQq
yYSAnn5CWoo6ni1+eil46cl27lwoecMCKKTaxTo+k43JDDZvyi9oCEmKEgUtRWlmevaPJALFin7+
dX0fQAI2rLG9FilKKr0/vgY/688mgqElsEg+l1s6Bw5CRPx28b0j6OlOBWJEj7wi5t6zODCNgh9V
kD/C1rWZHrqUvVv0MvJvVhXDNJL7jEKOQqYTukYv+kLll+DFUOcw0pOC6g8dFTbaMzYgIiml3n9i
AzDmMR2vQ/rzbv2HxIBCvKZUFnnoRS/t1p5fj+PhhDzUB0st4jih5BkvaIP6yMNmSYp0f5RsmfaK
5yn+oSTISYa37HTuZJyKQZdGVxZ6trnY50874c6a26t6mT98H9UuFvt2QkjhNYcYadUc8D8TqmA6
/mXdFWbEg224F2KJ7Fxdx9etfaYSou+wAkI0BMO2qzk2A2mRoy8BCdk1SYduI8Q799eGG/IKAOLx
v2ZEaEynLBxytuD+o0s9qF/p27pXxyUZSxz16wCXZoekSsMp9vI+M3+CtbzdJrjHgB2TxAImW8zM
jBI/YELDXry2hhNzamBXoLfvilhS2OW5WFyJY5T+Ezk4xOCovA8jR/1k221PQKfbdxHU5KMYd8iT
ake0DOFucLYL9V6EU8ykci8U+JElSY916gmL8/+V17IIN3pJCpzVxBVXY0MswxJepU7pW9+LhLpF
g09cz5Z4C35Pqgb6QWciyLqSNkXADcUZa/kqAzVzfMdB9myGMetK4xaqYFZw+5qNnHM1BQKy5ANA
Jhgw1nEfNPJpTAvwqro4Zr1MvIeO4UUTCbk6ZL+D2kOYx2Yj66NnqG4Ee8Q6ALPWNf8LFcKBs+XL
TDmfZZNOnmUcbu4Jzg4Aj8jU98ckj+Z/KOFqUhbBNjfNg9DH04f+JLoiq47nsC4GJOrwaXGdvLMH
pNfidwI1s2oQwHsj9+u4B1a6SykEiC1doJZIw6BUkhKhNbvDjIdK6H6Z0w0g9FM5FQipHGbW/hfW
Ek0s/Obqb7dY7CPHBJiEkfgRduFzoHYSjj5mcKAOhuy5bsPNch5/g9TzV/12n6wHWTyr0kWgOwLR
pj9Yw7IOxXJgkGl/jl1Mq2QjviAPhmqz6fzANH4XyJrYw21ovrHS/1lxfCqw4zeKDiA2azUq3aPh
f+snoEzxTdB0X3A3fHe9NeWYm4UR2ZlVuwvvuM8OZvvHlgoQ8Ft8OO6T53JjbSEg79ttTL17MvQN
l58Stm72uQ2ppoX4p69+R8vrU+ReCG45VI3GlCIk9DtUmRv59+coQ0cL2TatMQa6jN0BJHKehxT0
A3DACKOwSWhiJCq1GY4tvV9TRV5jqPeumnr6ri26VU5C6i2HQh/o1rgS2HvUC887M6Y5FTQ7NXNJ
ZyVIqVL6FQzlpJ80PXxa8n3TKCqKWJhcgUHi9vvFwv+5DT1scGWSR/uE/2lxdF+JM4ksz+G8KzLQ
s1deMZtFn2+1skQNt5QCMcLxaJs2u3qubOPAhizgxFMJaqPAh/SzjXU3R7j6zGxOGmlpI1LZTFxg
trOd447A0PvlqB7ilUZ7UO8klgmTc3u3Di3z47ZKpJjFz/qGMMX1AXkub9y8lQV0bm/3wihmyXz3
cwWv+sf2kQgAnR7FIen9W2OGIZqBLeuZc63DKpYRlD7ozvrTDYS/OQ+iTqRevKDY60LcVM9qaTG4
Y5S9ZWdd+Mazk3PPf3NUBAMLUj67eLB/Y04zMzfWsdgiKL6JIgEs2tQa2oOcNWaWy946GXEYJdp6
B3krI+wSCoFqfIccLj8xDza/Hxr00/W3/gDMd7cxyIHKgivt4ZA0V8GTlVMndgg1v21ECxlj/sNX
x/YYNZbQW6rDRkI/7l9g9h7Y4AzX1oXqEUmtsliL0orMiMjNK6nhF1FrvlElwW8nbb3sOhCNX2R4
go6yrH8/1VPFaFu8YNbIF01jeCyXapVh0QiLBWRdnpPPsH9JdpTyLf8Qne9VHoBQOZNMcpW7rcgK
Rud/OoLaUmmIijq12O7Ur1VLtsLe1rz6ghXniYs4xhKaXcY8598Va/cq7cXqww5DE6iuU0Tp6NlE
EkAlXzMM79zilN++k1k7VGMPqbkxljsU/dlYcnpSn4z0S5tEGNC3ubGHhUgwmJOQcd1yoagmdhiN
Drs0uqoVQ/GVT9R9zLRkVlgnaOiCXQEkIebwjsLb7k9s7wvcVFu1nDnLXGZtBhq+et0/dpTKw3uN
GSli7FE0+UshAUMuWpKshEMw9YXYnR5GwP7O5Zqsil8WX1vWcH/AmsS14lFyywcpp1zrY+jqYELH
g7vbnnq9xsQb6j4ITw5hJB0Q7FFLqsqv+D1oM0gPWTqzWz6Jk7Ez4EyRfYpo81xWHVJzb7sBz0vk
EqBfGyQYhTEjroVs+At283/h92YxXlQzktEgInlrDzUEO6jtu5ZX98REe+JVkMFJcNWAPoL58aon
mysavATms9+tT/3oz+RWheDhfZ2SntYA/CAwOTv9/q+DJ7DulnvK/TYrmXlJ2uoms/DRMcxVfoZX
dWgG9BYWLrB3z1qZqWUoBuUvGnAzu8JokaSQivJSWsCVzJKJ4z+uisfPhm7+9Zne/jO9iFjFFz6e
zwyZn3r7N5vH1QtEoBIUq0kJccsjTzV847G4qYMQLmV/cxAnFN3flnm2LAGVeaUoza/wIFCGL9zN
sCYLEap+0FVIZYwkjtHzqAvv/FpLuX9XktPw+I658F9wKHyQgPtFleQ8sEuoAv/OfIurajJAWL5S
f31leyt+CZwOZsA4aaVl0sP5QYmoVg47j7XxTVzDFDN26hwamaxkPustLiT3jrntbUZZCPLJiLjb
fRTD7hzWsYw4PQO4/VDkaVQOBmK/4HcKNpgZmjyeXWiZDrxUlb13RJEkBvXtk4LeLB5V5qSOqbn1
iraR+VchnIQ8gWLSrFUODI9VvgpdZwqMzlXyIfv8pNqM7g9gHPCiahriH0cGlV6zmbWeDQo7ImbW
8T18jp/dghP6XoZXQcFRSgXPhDAdR2ZhZLCwMxiaCA5WlHn77vL8fMiMnnO4yTH5lzsBjNgDI3Lk
ko6AiITVuzSMH2IDVS/wGCzXN60KGpZ5UKs345xNYg5rznAolo6aj1Oh1cfEB07mGzcJtNLVsW/D
rViHdx1lzGQAxPH58KqvHUskswvXW0BjSRIAcABYLp4hs/+AY137tfIZK+hSNLvgnI9XWKzF81TR
f5o/1pIIx1nRJGrlgguwKkNT0m8/7B2qrEe5rqdAuTKpn/7GkPx8drJcwkDhl6pObtvWpSScG7n7
xFe7KEIE5hIlNDOvf9MFBnAuPGKfb+GWhMuI6JHo8F+bI/N000MHDL7JTvETPTGrqWwVN+cw8aCE
UAfuUv3rAZilRCAcG/+DbE5YeNKLgmjaKSUNRll1lMYFeJbHptoAvDmkFUl6DG8ml3mb16O/xrnZ
BJ0CIFzX+lRtcUpT7UqTMd55O1/BjYtvuTSCEkMTHM3jEQ530qJIsiYowYSbDdrYKbUsesxUZjjM
O1Lt3D9RrS+muOF7w9wkz3qKbn94RCKn4Rpa+GPdWrcarUXv/4VlxN+cEzQBbxcXHPCZpSN++Ag1
2ysFHZz/N25iWhMOF+1WMZodt0oYvfF+6QctXqWE1mH420yLPDohGIJD3ri1GodBTPppZjEzz5o5
SzWa8TYRufpogk5804Z79hrPRn0XLrKQpiMXRjCsj37jBEzNAjXWXrw2pPigfXEbcB78LDlLZf9Y
1fEm17OxMHV8Nx2YxscAzr5cfNKhIdp0liO2HTffDEPeDbt+iZyvOQHFx6nKdsQPr9297tO56yY3
uWuc6CnSfVA7imEWq8KNAAatBDDkzsw4SUMnPmWu4Jq9UoGEBIxWEeP+v4I6zA4POW7FPfIIN8Vh
ulRo6dp71dRhplCWl5t4MGLu40dWmnQMNil/2luJZd13iWi2NuYRr/L2xiZc+/KsMzvDcPEN9EVn
CzMtbOxTuKIjtjBIu13i28uHbVpZ5RVYYCJhYgDEdYVH73GHTXi51qv4lFWTfXsbT40BNsQ41vRJ
KBqM8S7MGcz8uTRjkOzblaFbUcmo3DFnbdK1JMUmEXAJjbcG2zOsPYQmd4trJ/J/U5xuRRe1UCRP
H1xli+ZXeCcvDT58M0ob4Asfh8VOUoMOr57/rJrGMSodYtreR6crNKK4KJTZgOlNLtf9qDhWwdP/
o3iT7Mscc2x9AQoK/3YL7JRU3cZTO6L9cOvVqfhgk5q5CbVetOZNkeVu27yG9QwVwjSPYXI4qtMI
9TfMxm5gdT2LCpW1V5o3WZgPQcEjhmUP+wRaRunrsds+qlWy/gYND/TRhEH3C3T/n/EkyLcaH/Kw
XmF8JGQdys223ZI816dIFuKJ9ZUCTKMGK9+Yif462BXd+ZGEToR9NH0CzR9hUHk4/hZBgLVTiMZ9
dwLSL2E33myYku9hOERFPPhifQL9u1pwmG1ur//ZlECejXdnzeZBm0rLLPc5soCuVxAHCFH3Omn+
f8/gD59uUdDwBe67aI0DKyMPJdg6n0InOrAWjvNuO3haFziQzHJr/jujY0MozMPZ0LZPp2sUdCVI
TUVdR0tkxAjsYuwh3MnjBGIJ3xdsG5L0zTLI86UuxpPSAmADVo8S1grHlXOaFDkpVQ+JL58SZCCY
oId8DwITucqJVrhvld3megv7H7P+ly5IYPf0HtkzQGTl8RjoVsYtcJBSVMsSE2RBXUmHz8K8Ibd3
UgxlN9bqYEBflAJ6uo++v/c1Os7vV9uaMcES77GxDguYcp5aPl1mTZLDtwouQv2BkZ/Rvszwin55
ZhHWmdpXdoVIfy87xVuMVTJJrKoPyyVgDP8QbVekzTW5Y7lYwmuzJZdEfvo1UFSuBXynom2GJ1Zu
rt+NytlzoilxYU15+DkFO4xL0s4PRSn82kS3Egvvvub1zgCVPnTa4+I0MOGk5mR0bUV/vPIsfjCs
lAxtWqYxjgOUyg49EO8DeeZCFEiTXlpROxWuQqXneJ+jTY8q+dsQxb3bMlNKq0TInScTE4bxMcGh
ARea1B6QkSgv20ZrUMfOM2I3dL4xjGnwmVMgyOhbs0ICsWTysdA7QJGKw68jSVAQmInastyBDg7T
xU1badbfnpxWvfzL8iPAJ+Miwea+/ziO1OuRAC7xwF7UCZ2WeA3zoL3ZYmZz1KEJ4kLunq89fNwg
+wv6rZZ8Sm6o6FY1ang3J0ATlBf9Oqz1PpMsN0PPvmgPdsKYoGeMDTLUle8Nain9HaL/bdA9RDja
vBZnaXB5LNhwmEM/1Aez5G2taJG/hBwHPOI8g0t76TxoXrVs5wxnI2fZrQDLxoPSQvrbvR+kVla8
pvuiUrgjVePb3hZCy4OsVDYeRv9s0BRc/uuJ/Y0fuhO7BZjZkDcAyadijaZPVvnmBIWLfkoQkMpd
7WEwjhCtEzXYOqTRyp3DxJuW4Ezle55LwHimdDZJJdZZ9Tkrr1zvhSg0x0CNYEqywhafrGSckc6l
hs+mOpKSLPC2iYrp1c0FFxN4/X4S947dtEcP+9RA3gpYbnFI2I5iBl/NlubTteXGx+BNou5DMPnv
+0msUI+D9iFsDdyCXrIqRKScWx2n+O48LBUKY3LJRaBZNfeD2ZhqhR3M3YqAZ8PHehRDz5tIBylY
p2dZsqpoM4p2ZRQv0zDV+UNG/yLFRoGk9504SY/5pG7M770lgoESj2QAfAUpdt774O0c247cTEv6
ZwsyIwgRQUygsP6ATuYx0NJeDLqlHRSngV0T4kUwM4iGIGYdPMD31QXfF2qIhw/1apzw6iBBSgOE
Ac+5x/j0osgQY7nAvVeiXq7wGGWhEMxGKtXUEVyddrgmgvg8ly6XUVDa+Ea2DyFpSHexjlH5R2SB
LHtTheC8TXGX94XHR34hBI8c38EQ7G6KyFjdFO04zYHoeE1bNZA0DznuJPV5FPQOdS3b9qQTZWBo
49zf0AqsUX9GBPz6T3YhqXXCqBywnHUbuh2v7IFlBXEj07vz2iNFu7nABiZkJMjR6v+7oBM8IuRC
qymBS1EbnCRT+eD6ZDwH7UjivHDp5Dt01FkdFuPkPTaF5jXj/RRyNyvqm66NcvuVvtboyS7Rcm6/
exDc008/WqZ4HxVy62/n6WY9zy0h8R4INNcHM8bpPpjTzfbJafNfN/BZwAbRSL6NFxUMkUYczvb2
mmyPRACZRKukeOvkmj6IIfzZzTpBH3yEBVaKhvt21+l13wJ08HBU3QwEri6/GEndKC+1loJTLc6j
USiDNhQ/ealxq/wdAovhnHtwS3SOWsYYDl9bQs71RKHlKm1LJj2M+J7ROQSyTw8AEEeYQ58RUGiT
tng7uVYgn9ROe0T3gk2ZTyQiBFSZzrrKCocFdlOVoEOIZsLF4Q1OmTXJoWv3EUGda0m9XaCqId6l
wPyaZFIzJMjckO2Rmt1iT7+YQt8m8Rr42wiFUpvMsJIByFR8e7N/R1SEmyfzVFu2ybpQ0vILt/k9
6U7G8ZdGrNzXE4vaSV6Us4QhVyAvGqhgbs1CfFT9kSwwKNphh/n6TPyAM4SvOJS8suiHGobK/T3c
q6gQJYpmqEgK03Nt0eCRxEqndaJcWrFO+PlmLyr1ZUN6jg1OJdqTtcD7/LdtEa4cKe3gpehuL7Jn
50mZkoMoff9GSwKAjKH/y83+XV2OXy7j+kQa6uYdQtZdJkSPSIXdsbLANlYAh6tVdArQ97x8rckS
gNy8lb5e6OBOu/8Frh2F11k0HA0zpJfhQgN1/4izIOe8lMiMhGqxvylm8gPVZ8t+BNiw++qNNRBT
7rvyajSswDDKd94Qo1bfRGXxTnGYwG7W07acgDgIZOAqyc0yNYP58R3IIXHPOZ9ZeMi+n9OXCjlG
Tt5UGoBmaL4HunSwAP8FnRF/Vt5KsKr8AM3X0g6kUcmmaZi9T4CoXIrO4YgAttJVqN/MaCRGCvdF
41RNhir08HGOqGYyT5zSLPKpiTnmb4lnbF/3QHOuvU20/ak9DL4RFxz1b3GarHjFkaWFU2dIG4et
xIx61jm5pOnjj+7ZxuSI/6/VZj2kV2wW5IvPiMlJO3ydD88X7Kb6rQAz4eHOiR7iBYCmttwIgSCD
7vH/8VivJIys1JIkBaDROdoCoxmwy3VtY1IJxx+7trQlV1YsjIzkn2AuYFXYuPb+wV931qYT2M8I
5VZj5D7xCEoK74RZ0iDW2ya/k6TcGMDWohL784RS3zOlEbXcBa8pkjiRoB6RU7yK1x42PLLydExa
5N1tS9/3Go5DBVpD5MBmBf4Ggbny44iXAOfY1zwukO5D/qIldf8+T+iFCF14yWA8Ceyq/962yWL2
w9Gyk4//JIO9OBXwN8fH51ti1VCzOpnRbbXTqXERBvPMQKQq5cL9lFhWGWExAtKr2Qly1d9QeRdx
kP+3Bbr2DwEPM5yMpzCFgdPfRBnHt/g2b3KLYWoyNncW6qIPLg8vYetW/emRa5DrSbp2gpZZBJT3
PUnokwcpuqlv1qw2gZqvtOMBKZOTy3rEvVZI19qxET1e5p65zyYQ8fA+WEP7c1Hv9JMJ603yh4zJ
28iHF/tTy0N4Pm8/4n1xtKaUX2bcp+ep0AuWQHtmlFiLTF1xPW8lqbuOgDNjFChZUisZnHLzQgqE
j/zAd7EzwN3gPhh/BEsk/lojbF6T++NGV41FxytsqTXEksTBRiqqgNKJz8OosXoO/wIawRD//VSr
3LipBqlmQdon/2YTztLTqITsBoGxC5t/EGCgMYd4WLWIKix8wCX6jKase/estCijRMAwW2QWLbjN
zqphvtRM/HQTIwGfJRR9yme1GwvSRydmnAeFTpSmJvBKOUWJ9Q3hjCDEfEYW6vRv3Rsqr0OS2ipC
SmuWxIYYdzc4F1wp8JkItHVnkFXQ46JW2nVOAoRRsugydAeFHwi/Ia6q0B79/f6/RIdvvEA7sDlc
ND5xqDIlPFk4lgrT+pfw2rJB1GAfvi+qBztpRs50LFXMdXFV/9IRPZuWmUsdU+FJQKZ9xHd3Y+AN
MNIn1a01y8t+ILAJOlLP3BfqnH2hvIno6TsXmB3O9yIyH7wY93Kk1v7CtZbRQbXAnM1QEG2T+lCY
EGV+I2cAyZkIQhCtyfBYznE81vddFP+HJt1FAAHJFFKnfroAbDyeH3k+N1g+R3Wxo0vQJ0JB1LIW
JVcZrQXU+tWWLm+TbDYeaW9PCCWpjhzD673Yzjlr/RHjIAQArNzUzbOAatuUjdhO3nLfTWz7DOfJ
LK8UaFKGiVs2fXbSch+FWR+yMtDvepzQ1FskYv6hXG0e20gSrnX8sQHa1rmbT8wYT7+xG6D3PhLV
OyISP87dF3eu/GAuIN74WZ4CoH+7Qy2g22aNHlZzCXnJ/wlupkHqJc0c1dlGekuQ3/7sYo5F55CS
x4f+sglrgh42atrh6U8yxaeEleQvwPEri9d7NwzP9fp+kFVkDWn/5ca7JvPxi3UzTFLv26UdVadW
XqScbHxSj90Mlycu6EnTzyiWJ2o5BmUr2WlT3A1NhzVY4NRbu6nWL5GaJQ1IKRSikTqh2yLja47U
EkWTUTRHTubXJEZNi3dmbQuhQzOksTCBR2wt+dnvJAb2e0BF0AZGK6yFmMl3Jizo+8G2mP/eLG9/
2MWAnNBSla9LMYOL0fe7ZlCIOsUFRzZPCqqCyli5jH8kjKJjOu/CYOi97cN4As5EnCydF1XyxJtV
5TNOqA3wC7jW8ndMZyzoU8uBpYMGi5cXohcHVoYLrwl2gbcZvY6sxq/+ksO1rAaBSCGgrsfsjJ5b
YD5REQdlhpNsxN28z3OvTKn5DEqI7XK371FRz78GhzGArQ8OolIfjscvP/E/ALRn21ki/vxe0I1m
NDlhBSrYK09HbAUhcMq/tHEAIrcCJYSoNvUiZdFUf/xiQEMgk2ENsanybw7Wc49kdm+1Ha8cFj0U
PM6aTE4U2vfJ5XLzu7xY4/3bllCcIez6QiYOXbRjH9Te81Oj8IHSa0+AtBpfxF+zq/rzph7fSm2v
hdUYZki+aOon+gs3W6BTtrM7WoCA245HuKxHI08SBrecCY4MmYMC11Og5XsOiIhygw7+NahJXuHF
CXdjVjPL0J68pmw7hFbgOJNPdm0qpzIbhSmInFq/jG/XIDYFtNT1VxcGn7x1U2+rFd9BCvZhEoHt
vPkKVhws4CT3gnMvaeRoc0qFQlcIna3ll+LsioSQcSkBbMeyU8MkRQQ6Z7rq2qvXGp46Znnc6+64
WwH+i5yUUYNv+vrE4pJOCf4oxX8PeRu6MVCeKaBDLY59SjfaYJ6EC81u5ZlnppiAZT1NK1guS/AF
eoEKxyahBItK6UdeJ9pbskA5LT4FDj2GAIi2ESvDwWgtfCsDAhdn9tQszxG+D8UiPElytosLEP3C
TeQCfy7l1+Bpf5DxZkd3WC74J1q1AsUoydhCboK1ERqHFybBLt9f/Ww8ISLqGYn4U3S2nsau4YwQ
u35UM/AKXpNv+3QfJorzLWFUcVqir5roWs8iRqb2uBcAONaMsIUeHnWtDD01oMtJKfCjcxgyAzb3
j+xE3u8JhmAqINk/Z+aweeCNVH7Nj4TN7czAKr/zEs/AIVQOrP6ALg4rX5BHhOto+lURyjzGjBA3
gBTkH+8HLt38U0tsWbwcxqTSVJM32RFRts2CoEh7K0Nemz6idG2wa19dQU3HW4c396QiY9hrvSJ8
mhLdWcI88fjFnazEM2uv8nIKnbaQo70ynEF+M4ZlIv3XX1EvoI4oIGBnjnWcex2OTiBCEfkmnBY0
yuhhZpNieuVbmLizfoDCEklnC+ZIyC6G9Zo6gaf88sqqq4au+UGbeDyjh0EjqLJfRz7onjwD97Aa
vQP6Nwf6fS+IVE/mzkKVLnt3X/Of8qK6P0uFCYx70LCQOvOZllczhBfdfcOmZ4wwKM9TMzC/jhjI
WNRjv22WPypA6bfCizH6IEaoMzG3JXvqirWUZ4+r8oxUSsTco/SYJjOmvMM3IvpNcy0+CE2ocwMa
MEJNHZiQwRUYAEuIqDc0fGm5X+Mn/vRa2jEfKeBn/RdIjZtl64xhIBn87K4Hwcc/BxNZE1EEhzQF
UYYx+nyvziJNwG6IEVC4eWrdbR9DqHKBCgWNElyaBmUv/O/FzzBgFAt7JtTg2sJAYfsvl5x3TcbG
NbNhRXedewze8BMnU0JcV9PK+VQS3Knw5F7z2j32ki+cg+vNz5p/zfKjF8C4PkhQz2kY54vnHZyt
6iE4uNEURbkrwkY+8a3HeKsD9EdFef3rILEl4C7vkjj2xqqIwhpgsOabeGGRHp4nBKzQY6FLqDRC
uYQgJjrj7WJG7HLhApnRrHzi455h08b8C2SQAj5erf4mQOG0tE1xV8Uja9IFmxHuCLFFdGrNmz5j
fexPkBTxfmhY3y8E731erfW65BOSP8LIGkw5Ou6l2DH2tvl5anEJU6AVuS95OtZfzextUin/TjDv
/Pu4GjS3LgFaKJNJGfwijlR3BM+3fVLvcEQ8cMLQTv+ifHq7BSp/kkWtlBeJeuwkf5zKISk65DUx
x8go1fa5bRe+bFAeLxZnoNEtAW4cLDwMCuTYbVF+29zkZMn19a8oJHh+FTnIJMfdaxlsRpkOTihU
1FZ1P9oqSUB2T9UsTZDH9H7tEwUurU39a4Cyfen4WarV/2hm5qaVDDR82Icr4XS/g+YXBwR/+32R
gCV8q1yJSMdur9jMyqOrY2FP2bwu+mtQqEse94rqzSUCSQoJnr5DFLK8oL97/zyGpanF9Imwg97Q
r3wh4yNg3bdEULWPSkGPMZRLzJ7oyPfrqBJyV9X7L5sqntmhHtVDFEeghMahhsCCdJNhQ1yP+h1E
wVqM2ewI93LF28KsrfKCQ3+5/DED8vpOcKZU7Pq+yD9Z7rci0tIR5jor0VLoFmYWrr+cafiMaa/y
8ggGwtE6FwlBLv7de5+0BbIQiX78VctFmgjH9a6MEiI7jmt9lMIqLq0uweiOGGAuZj3PEedsdrL/
44qiogyTNS+JT00u+xO4i7/bNIXvruLrcrFO9Q0Sk7iYViYzF0nBoL4F5uDSQ67XoHCNF+1U2na5
cWChjCMG5JYIJ3B2NIVmLVemJI5SsKcAn181/NOvA2fHR1GcUBDu6SWOPCg/Le2xW7xuONQdX4EN
g0Qw+Q+jz6AxWVIeLAMZ1+/ZzMDVEuku/ckDMM4TLLwJtS/JUjzXcRrX2fouHVPgfPW2lEIgmS2t
XQDjjH9rOWUGHK8h13sWQrGPs+4QCbZ5gggfdxWJEis53Lk2nSidsjA16gygLSJlLUWgV1tAbi0P
ey/fdkpcw5E5Oi75zUQWuMhaLZjLGy3u0UcwPWbQPAwMh9/yOD5WEsoav0SwcsTe70avUsRId60o
HHMioEe+3yLW92LFBsrzuqHxWoJXXSsp8GyQ26fXg+KDFtRfq8+L6Qg4PVMUIY7oYpsS4X42hmfJ
SKHqWRphd/rUJ8kKmIaPxeEZbb5H7+rgSfkkJsKfbQQtxWae/eTqlU4if0ZuEyXcgnvm3R6MndJf
gmT6VnknaLW2B9XkvluoVlfEG3UmbRvQYbR2RSMRG+0ewXhp4DpxoEtZwi28NqY1uZDWQcZd7k0M
I/cYWGKc7/VM0zUwvk8RfnHjHGZhNISDp0173RwZ/YOy/AkplqhGeXA4unEILd6WoSPMQ1LxMDB8
0tjPI7Rk7TbQ2bLLCXSAoe3JfRQ8Pr3GUluydyVTwzkZzvAfZoqUl8Z77XIlAbWdAwwP+oahC7Ao
IXmziOmwBkC3XEvkhHAcjKYWkYIhPL5Z7s2sLMQSqQewCSLrRq2KaSHwNDlWeCr6qVXVjx7synhk
z8btkOliSqw2grATOoxnoDExKHTseTOTUzqJAtWhrGJQ+mXCUmihNNhMlMEeVKpkpYdei9Glwwu6
GWtJuC8t1fjFuIJxB6El0A9ysuaPZc8Hllkie43ebq9a9drtXZOzFHt+tEuGTJk9Bj4ero9VReuL
dkIZg/GdvEB54PtzDQfsgDxfNUbH2gzA89Cto4QO48jtnuvEzaFmD2UVEDYBiZhTLOOjp/HpSWx1
w0g+3GAQLvAfTYZuykl/gp2SRq6gYcbXgS6OPKY7lETrA5fTZtW6xpDb6BBCKn57MaYhdahcxjJ/
cQJT8zYPT1cQ0P/F1tVdTCJtnsVE5qP4+doDSzhmBBQTnT0IQwVRAaK1kqulnfNXHd/2IRn96NrC
lzk+P67GNF7xMZ/Ync0su5VR7/eOZDaIUl7IBTGfPwageH2LfdNxC/0g2Fv0eCqTA/Rb7g+3PPfW
q3FX3OSvOPOhIegQYM/9jKIDh/WIj7YQkEXc66Wp4OhZwjUPRDErdE9IYr10imv0efBWCbz5qjRN
IRlh4q8VqyS3WmGpISIc7iuLPHbnj+wjgvZIb6RjVadqfFHMRxiVEXBP0RXpw8f8tbKxbJN0VTrN
KzNRDvTlqyKgBFW4S6Z9MBO0W+QDiwdJgIvtIadObtwGAesM1wB4U6PteQE/VqneqBpn8yoZKj2R
GKPfIYDQg1GQ5GuDkqrae/9NKlhOTOPXjgbHRJTy0YKyZEUH++ESN2u62HvKt+wzMNC4Zsc1jfU8
V1wux1UvBRGQ+xQlhD6gKjoleToDAqi7SzXhXJ26IgNANK0CR3/ozjEKYM+iEcuAnzyStJg240Ep
sf0nHWgcOwuAwAVf6Hf8kUkEJgDFrFQzbWqpOAkmMvhXtlJBXXrfL7bKp6WsrxmroriPNzcwf95C
bRENv56NN1m4oidw4tqbofID8A4VXl82iv3RP9aaGUsc26iUWqOVjzRsVnRKMnwQfvM7L3Ndsk5I
W/xZdF6xQ4MaMeyGDKf2lObthI/A+FYxx4f4KFfVt/UN+4RtgOd42d3bJiZIwZdsEIRXb10gn3qK
EgXyE22A11DSl+wJKPJpTPe6TfHYYmlb6gvldE1qa60gBPGKrwnJ4i2i0tZ3eWpqqSMxrpDd3XCB
6if5Hht7gq8xCYtCW0U27KOFElpLJLxWmhXafHf5OMOD52AMoNR76m32Vtu+xX2c+6FzSjWQDYhH
EBTQOlqmfT6nYKWIPprUbOv6KsrTAFIMUH1cdS5YFhUrcL31o4/W4RM5tsZs5Qu3jQpwg+f+hwvd
+2wgGDAGvSuDywL3Zzl4Pavjkemu0H1jAq6sruQ7kwAsKj5y73kY+iVKa+NbJkDPjYs9y5kSmEZ/
72XAdgIL4uTTRNvg7Kq24ZDmc5b84EZgHsH/Sd1ZohBgvkBHojh+3wvLQmqNu8aDTQPXzS4iwrP6
mW4VMgo392Tcwvi55tLL5uAFR+mxXw12EXJs/oxmaQ7ox8OUOVyO71+QPQhG6IrQvdGKH9Glr9XW
GOWWvCsqHWLx6lRUy0r3Vb61KiLWUAr9KLrbJzXXEGYkDs52tq+as+9VwzZOe677xXKOvhwSztW2
UZAytDHE0J7/IeilsLMyyZJFl9mj9buZ1nZszWbQuku60hgtuxIRUGvmXKDZIHKGD0bqKceBTihe
hbVgximp/QRPE8xldlzpcSh8f/nZNoA6yoTwhD6XGge1BLn+CxsFmLPGCmGsvSN5WUjyHiO6Bv22
czdQhUK/OJdy+pRsSMoknrl7zuHEpb47btHrKTGZExMpbVZBJ8ovot03MIlkvnFSRWDf8XvcQ9xV
ZgPzBL7ZSn+P7rNa51YKkJZKcBeW1O9mjtcwX1NDYO5dU7dg/lGVDC1UzHgDoUKL6qGOzh5QD3cG
imn4m1xfy/p1bMSxeJTphDNMmrvu6r3KBHO+tLCkdgR2/EE720nQ1byJ+LH576V+AlPL9Q2Ht1K/
U7UwrsScgEXfB/eBPh6I3CxftiNzles5hpEkyM7dezVkjUA91UMzRX62ZK0HEDaXUenq/LTnTywx
MTLg2by1kILiVBSpAbSkOxa3YkEeBtoUYXenaKQgtqRGU5ZU60kqZFfK6KSqCTZeWqIqgAGVbIev
NN7BdNZB5A9t7QXarEyDvciirhgLb84Gs1ue0dAUgB85lzgttEy1E6/accAc8ayqr9zPZTvsZJcb
0hAixZimT3W0lf386jdNxk65NVuM2v+UFUU7okJiMH8VSlHbNa2z3gaMx4VNfv12E5fm7wxoZfcP
2FvBKouFep77WlsrbDrFr1kSK8OQL9L0TtYApeUi2dyN38rO90kfwcVV92+T3ppyb+REr80Jk0sh
rCUYgI4M5WXh49TNqqgupkWkUQppfjTQJPrmYc3OnmQDvQiZaJUyacjbnUzFDjF22xn7bHhLcgo2
sTRP9heFs5xDJQEowfoPAC4gyjUArZfV0JM8SXVb+Vl8VMQkTuiLTlWab0ny0/JNwh30xj8faJmC
s5byWHEST8lwW8hJCaIpUtmjQPMDMSrNxNxMiB0CyfmnKWZ8cXSNdQvnWeKLl4uepzqZ4MUUDkU/
y/RYwueOmKqRpghZw4NYGcPMXxoRVsnf+2O62j3QQXLYw7YaJYS9qV4HK8eeRF4R2/mldTdwLLXK
zhw6QKbVdstyfSVeGNSmLdy7YQuLwoiR7WpepeWTbXlp0Wadg2rErHjlMZOjZUWgC0LNzC5OZXzo
7tEnnWi8uU68eQQo1W3kIYV/QtyqqekF22pf4Fl/HB5mt0ZGw+EJuGhGNW7P9S0NbiKCO9kiC8uU
PnMemPSPcz99+Jz9Hfw8+8L4XVQwCQ1ZyHv1fWJDhO175cwicDgV443uxdSYlTrCkmCjZLouQ1+R
lanspDXm0HpRqlq+GGLQ1P97aR/ECUM91F8V/3ppbAa5W28FEWnZA45sbhrcOMKo4QbNiKmkPSZf
VNzCbCdHnilzoiEslH2y248w31UUkhHVqsGiyzCG67pYRyNYZUr3GDqgK1w1AGiabgAGJ4Z8fPys
oDnmU9L00P3jsdrVl50p0EReciN7kfm4Rns+dR09V74s8uLxtCgY48gLmC+oS1O7qTrLltk/c0mu
/dlmfvs8sjI9ZXNP1Ccz9x/bIUSKaDUnABpn2F9kcZvTJkvs8bxqntwyd4qKoIUTLjyGX2+yoe1D
qBPLzpK9DX554MGMD+Ks1G6JOerEdVT74zRH9qQFQ2ogx3B08juFpSTH2J022tI/vLu/rmCFmz+T
v8+1E07tPfgalma5PACYBWcc6E2Sewj9zjLYlHGxRSKWAlYI/oSt4B553z6zLMEiXg/6Z8z5G5Ok
dZZr9ENwfkGFW8WljXUbyxAVVH5FnZhT7X4MTmqnvOT1s/cHPh9H5zNW1iFr6HceSHVm3AKM77RY
nFtX4UTq895cRao2Mu0NpZ9CbtH93Sm0XATrxYjbPxqj4VEnMoKN1NUveWCA+TXeo2/B54GxOOro
AziTf+KdzLI7UnVy2Gf6sSIDlaXhk1a3vMmXMG0zB3ygTHPobUmmLrn7p9FdX2IfzBvPotePWbfG
xJQbjwKKC9DSjNDVfHLcOnP0SSQ2DV4YRbmmZ0IzbBiaKbgtwBnvbdcV/A8qkenqH6cbRVMk9uhs
oUFbwpDALMRAuKdspQ1bEDIkWs8O0O2cz4P6y4rBOzxfb/dTNqFdiNWJq7SvfFoWIotkDkj2OCTU
UTBU8s2oll++qKGltOceX/H9vmn5zrT9c14Ky1bJ8gWxjh4o0ZnJI/apjQNIwoHY28ORWI+K9Apr
gvwvhVnsRP7ryKDVohSwJvJynbp126lQ/PtLvjxqJpykTWei+VC7DQAPV39BtPBlNeg3OvCWGcy7
1acpAv2xQBAEzl5FHdFHpJ2Kf6NvKw4FDNZwNgTCatrwOfETwwskNJjEzByE2qppe+8QgN8uXJ7e
xvwhkoRtFpNhtcXmhJaCdEOVfSQ7u6wLQUQ7JBmEdZBqiFhwcLXm2CzmJu2J0r6Y4G7h0YlYwtjR
Ae22s+hsbKpD2Idt8rEyuBASwCGf9Nip0g2MHfE4JzU62fjRGqMLBHu3DDqmXbyn8MWMxRode1Ht
/lhcD4g8y/MOL6wEDDWP+sDrNSzIz9RlMMJSSpK5Qsaf+CiGrsHtQhVG7QqnZTaUZyg1Qaxyq3nz
GytoY7kdPj0IsT36R6Jlp3ljLWo/ONsiD/UeRFuR0X1lWgZ61Gm149627rYasvyJR25Pmd+EIGJi
PRUrOr34M9uNNQpirCR37g3y4LVxEFZGwrhJduC+O+VegXPSLZXT+syiyZJz9qkDsIKTn5HtUPqJ
8M8pQPTp8K16yAr1fyA/uWm2GvMvY04eIR+1F8MNIFpEuxIgG0y6E9voC/XSyJOFz0y+FcSch2gj
/gHlTw1G+qaWAC9SU2/dgpN34L1E2+ISo4WGgpHSl9BHUAu2tPX2Ynr7Xunz4xvDooBdgxpHNt9I
G4OYl+xMte+X05A6cVtW4zm/EjPhtGlpznfmYcZze29zKroJ9trB5P6r/ItzO6vkoTjagGJVlUrh
FDh/SSzGaHxc7Cl2nXWrP1QI1Jgg5lFPsFMddAdSUcUaabY2IUZgZI8a0zYojfE95rU4fdz621XA
9h6iJ6WNfQzP1JVUSc40kRJbMiP6ZIb7fOnCyNjhuyAmi6fTpELy1JLt/+OvqFxIp6PgEhiD/4AH
wMera5k23mvasZ5PPPH3EU95amhF53CX8uDScXQd7zK67nQU3MAs1C2ufUwvtY6HbXJQ67t9YbuK
pJPo6t/ID9vCQdO9iKUq+k8AqdAa1CEblBu7OiRIuukV7FqwwN87WDEzm81oHqPZh+uSGc/A9MCP
mPqyk27MojTKm8K2foihSRpqPri3JoQt/WEyrtdFroNq7vkUywggFwJrVsHp4zFxBFkK4ANQztNz
ITQI+Hds2ugf7K66LL3MiR9SIwITn5ycO91id9nP0kz+iDb5KmKV8sW2c5HJLUh+15s9m2KTbnBX
gjC0peJeYMcORKymhwtBoDjU2HOCW5RjYyPRpw3gbo7nHD1wKPeVsfNa9WtzbeLA9GW3sL/WBCC9
gdQUjJEtWUSyBEvNvKeVH28m72/ljkmBywLwm5GT7MSUsrNxoeVpXOum1T661HyIf9EhTsyAv1ca
OoGTBg6Z5O2txQhf/zbODgupC6xt8DYjDRVZLOC8ktB0VjNYtscag/xpCW3mc+U+0iMdqFeLh3Zi
DtWQzjXZifGSyMPVCnsx6ZMflyl4I4zbRU4pk2zoVFurEFkusbzEEoeGto8Hs/SJ7U9Os8TVZOOC
0Nb/GEf+Ywt8ytLdi3jz2NAqlY4hpgFej+JPa0D3Euavz6NPYN0Nl80mSGG8Sf4/OP5P18L0tRCK
tGaItYfOlPWBJB/1WU5DbSEEbdXQTbf43Q1hGBh06jdE2xDojQUWVPOS2q0Zeky7hw/uTVdyN0yF
zPx5VOwi8cRKg7KX+xFMsv9VoxTzEWqjMXMsunWxUXEfw7kkhBEqrUgJoma/joG8REh0vwEUtTbU
zw1a+hyZuWSEQ0Y+uqzl+uC1Td95V+UWgTj1QOBMev/S60BogISD+vZ9v2m0EwXhTngo796z2+RS
qA6dxrTHcXgxRousDHVG3xQhFu1DvjCAGhZmR4pOg2Z4nppTt0SuzL54jjN4mqfdprO8nGwpM77a
sYhfMVSt323LUZj/QDISLdJW5e4mN1DxmdJDEjdIC8gv7ooMtYDzP//Fubh50GO444U29V1P8JL1
gtogaqj+/8ttHElmy9tWIkjen8/UBjvAfrz1KPqvkREltUIP1tbAF1RvMS4sjNXzkr7vRG5FbGIa
zEt3rTpifAkWOM5wOLBpWELMOnqMQSh8vDY5OFGUzq6XG8GvF5B+MB7KIJ8tfdj9/wH6mnQtAe8y
TNuurO07h6VptZHeOC9DO3dely1VImMQ800JyTnsZoEZPKg1t87lUmVfrXdRKwNjdnazikEcnjbo
5Sdrnzsrv2OIQr+eu5b30WsBYM4yHnVveWd+/UUFf0SXYxr+gwiVUfGgT2w27ZZPOBjZZVOIrgAL
5la2rd2HXf+s3YeOH1Hqdi3jAHlzx6SeSmpUIzvmlLiC2HoPdUxdwxTB0YPzOgDu0PQUEiu/rTfw
lrdCCKAkE/f9PA381CqXFEn0UHOKobdhPmu+WpM3sY+9iidvRxT3uAugSfjbTcOwgHIPrvKnni1c
sS++tJn8+JgSqunbpyFR7DVBF1DD75Oo6pVEcumT1thzjs3RDh/1MHew5L6EV3QmNuFhIhNKmnXr
35yhB2L0eUina6ErOyifXrdLvTdmMFRNOO3IYyJLVXdfSqHkbSFAcJTxRJx7ut4oeRheYXrK4QEF
NwT2KgSmtnyAOAjpDdVI6WDWT1Pg22AOmec8fsCgYZjTUwW1dz6XG1j9UB7jQReGbR1tyXu4Ael7
FHhauU31kEii0Lb5TLyyMzLqu9I0JWSaf/4QoSdsvwPWu0gtGBkZN8S3has91O0mQXCR7vtcddtq
xWM8Bne0MvZhO6zcvKrTJ0C5/7IwjVO1DMl4LgcnCOY9jqNKlpqyD4JUnUZ58G+Nw7ZoDV40fduD
gW56W5651RrRLkg0VGKHwVmGEiaHrL2Dzbr+G5pbvSulxZRumq+Jkxu7A+YOqzajcpzdmcIyeveU
rMQYzV5Ei+7JO1bZjf2S+zh8gALMnV6uNUV9/owKxGjioYl+DQcNauFkzvAlA3zmzrixAihk5K9j
T4GtbJYYPKy9sBZ4HgtttPcriPDeCF7BDTtR4WKd6AEJjDnlLI6FIhYculWRyimaJEj1O4bxZax/
w2Pda7WVkuqCTmBNSnN1sFEf8ALf0s/knapmGFy3fAl9oFNr0pHAGk9HkXd4soc7F9E5RCbrqk6L
6G8WdLWqFL9A+p5zTyjZBF1u3oZRIMYhUiZ3DQzJRawDB9Va/TMVIosK5+If2EGQZVb7+WMyYtjm
Rf0lTT4WufTd/dh55DZAfnvNxHsr3XsGZTtz/Mex3s7cD8C5iXe1KqJIENBYedf/sDVxdAvo4rVV
2n7ZjTP4i3gQHNH0v6by/8ggiVNwVKvEH+u8f5P/Z6Ek75HDMjz224wAkH+NQPpti9kck4yGV3Ye
jG0OipHD15k7lzj30HzPcGFORCjOIw6ifsGbMWEKkw84pTvFnw57NvlZ0oUFiDlscw1XhdtOwDID
JXF/pvFNkSoG0LMoUJZXq74rteGxjPGZtPQPcBGC+7ZN+3ybYR/H9v/lEfUJijC9S/LRk8VQqPhg
WtvWY4yM+zH5eQdm7ainT0KB7HbM5lgCiGoYSwpq0Gi24XJ1+vCGq1eWVj8DP3Hb5H7C1InPPJSf
lGR19nmnzTvSrMmHQzNNoTfz8pyeqyxmbwXgeewMmepaqZkluFnrrqbI0X21rUsrJwmcVPWKlx6v
t2aZ0TadF7tDNPSQrglYku7wqF89MheMtCbe663dCggeNPGYdh8/C+FcGHMhdCny3XjxnrBjSZQN
omeR6EYyC2o6tQqxNLLOXcDAb8Qi8YiU7+UZ/m+sHivd35tJJuesX40Poepn5KCf8JDy6FwJRJuv
wg2i5j03r4hNoJYyfh3KoYTp/oTlS1TTLErzptM+7BsLiHmyfddwxw0MFmzIIJPejj/ZMfYwjhp9
u9qqoyB3HFqBXRZBYiOv+N7dK0S1kRYeWm69KF/EaoSQ9vH7Jry7dxKL0ZY27wWJu8CEOgN+zxxM
/gs0yYId+idPJAqP/Zi0/TfhcKTHqtfBPLq9acdbOOdOGu08uS6vzhvw9K7yd1NFIjHL82ncL3Wf
/X1ODANOWNsUbGmE2tl4tIqTK2Wa3oaVOVwb1XQ27OgdxP8DU1Ua+coucyOcetdphyoBDFPk3ftF
7KTXX80ZQH9nweHvOEz1jxlre+o+C8ZLGOW8bzLkyQ8Rc8OU8g/k3kEz3fuYbW6ZHDnY6Hu3TOdc
cJ8iDxmOrGGYBnluiq0PKIwLAZaFyerNiI7Wvoep/3vO3ucY8oPIg/owkYDBfx8yi9+w27JGExE4
r+h0x/VWiQFLs4pxJUnB5s8hFzzx6S0atEl/LXF6qalTnlTCF4rcKGeoDdSpl7kKymGx4b712ky5
PGhenubzAdqGrlDR9+yiuF8iZs6xnijyoJaHGgBVw4A6X7xzCZqqOIsfp5dRlFk/YcWY6lzLFX+A
ZVaEFSO/G6/jxaWzoEDWOHMo/89XQiJHzIciLyM39EazvPE8/FquoWv6IoUddDiSqEgv2G3M7MDa
tSYR4MDoDAwqes3qV2cuTGjlU/iOsVPnY+6ohfnqA7ZwlBRsLJCg15OIxvpDNlH/VTaQMp6louW4
3mokhwes1mG1mG69PPwhinOLnuwfsfp9RAHWUhF9f2HixXkeYTqBBHdpIrjO5XuSGMayQEhsXA/r
RJqHNQEjhqs7JwZ0ZbuCUftA9v/roM93shxe1c0gPT1nOJ2vfdLrXQP1YNsL/kMLr526lqrqtE9J
CoKzi53D0GKuznkOPC22aGWCkvs7VgURyOf8TkLz1dHJ0BWPBJ9yUusoPmsubkIYcKDCvGLEu1Rj
CyoUeHnwX86zcTy+0ojBaiMxlv4MnR8Lio2VWf9Ooeeb4agN2XCxkr7o7BqSdwzDOUUoIgCTSkgs
pybIbtlIRMlBD4++le7kCLOn55H7q84kgFBJGnc5wNOCBSO5hwF04K6hjdODagJUCv2GLTuE/gA9
RrGclj4NVdk4UfxtEXJ10HPpWtiuDtimL/U+T8woDFGKPVt8QyJTXpYDFVKLIP7Zea9W1joCPt1x
O6T9GBAvBPdI5Wxf8yPMltGFQpiPHCvJRdfk1MkB5jqjCsSWyNxHfzB+52JGdbuvvm1GS/VrWDI6
DI1sgf5pj0eBywf2bHsd025PHrCgNMFpJPJ4y5zC8FsvUE2UDqp3DT5w0vEMMe8l3r57+pTWIUoL
5TyD1E0yik25pY5yVogUjtt9vUSSgZkNvl5ZCYxrC+2IX8JdyA6NOov7JHetqZFRPipfHM1XpY+f
DclOSeyG8xTLiKInKBBksZUITX4UCMfTH1XQf9TTdpi2g2CGikS8ra49PqHKzX5EaEHawvvEXlOs
Xt+nLzsrwlMttnYy9I0o5akOg4a9wBLt5/CbTAO+1AtwTC7Ic2SJjH6U0wbeblz4HbDJrZ2vMh68
xLaPlPwvbxUC+6pn80GFpRSEMUUgrDzNAA8Ca+liXkTdxQFOSYOYwXNmvHjNu5qgbPTWzSkM1bpU
qUJl4rtLqofOdizof4QmIFneCqHuNomu6/X3yfwW/qZKqUi0Q4HiFKdqU7oM4yw/OlpOtbuKAftr
PdTpoZB/QysUh5L5q1xrTSB1Rvqk20jgWwafklvMSJTaqYqlrtfBe8IBls2Voe6rWYw6ZKWzdqWI
nbH5pm9RSCXuaNNuJ35HXZHeAT4Fx6nYQhplcj8J0CrQFbQ5uRvSP7vcpLGzSd/UIS2GhVAB1+oO
zBRvwhRNXcAwS9qDri1aeD6G5PZ7S5+xAnFA3hw+vzsMWuZn8y3WtV7/P9hqyr/iivNYQNjahHMI
q9cPZ4KyejYeyA7GlX/Fvluzw8SQCFlo47fjxV9Vct3yZg3Mdo6wIYlLXp+p3uJBPlY5HFlypkyc
aiXZ76D49qqJoh/Vup1h8kGo9dAF2k13UOr27W7Q7HkSSPAdXVtAFiKpMxNs3sBpaO1bZ2JX1fys
IqtpXdeXzFnIg9BeKt2D1ODmnGmLJdc34jyZHtEKtTX3sf7PELMbe/Yv+v9TuQv6qZPHLEtLxuN5
oq9xx8yTYg5Bcr0qFtGXNTbYUXQddWhiiakGt8bPXPBj8bhQ0Fb5vZFximpEnz/BSHmia/l3fyT9
WFb7KUNraBkzaojtihVZXjbzjnMVuxSxs1QctAvts9Xrleteq83SF7szuW+D2oDSJ4aJ5PkTOUDd
e9S9nPFWzNSDJg2j2AQI8Rt5Ijr15DEnF222lUlK9lN7gNHJGG919OjSZMf4UzmrANkJFUu5svd5
KZ6AKVS0QCPmVzLAnfeMzUtRycxymlegSLRHnr2SFe2FjqNymHxpUuOmcb9zfL54/UOvXkGqwHEt
duF244jQrkKUs2KGt8JJVqwnkofiJP4vN7HLNdwMGiDXFdfeu8cXKW9oaYUIDGFj9JsN3Rjj6/7W
tHAZRkMJh7DypzqL2mv9iA5a+3omfUTr5yj2I4auB9PZpzD+yX3MsR9Jev2Gxd5lA/fJpgAE9igg
0XGZhGvfsCLiYO6BWAMAhM0KMlHR/9DKFyZsEK7LAQZ0JXREH4yyCwBAcxbFVMawRY0eH5s8ZRnf
0+tlmc9JQumgNO9Q7veOg+rDYu8woqc2Cud0sHyiCCquc636CpnMNE2qim8yBxF3Q22kMGiP0VmF
1mSkxsV2bzY7mZ6J9oyAuAaWAtVOxSi97vWLM3Z026QPWccTDwnRAZ011Gbki5onmdkBQW56sZjW
seMktlvw5eA9JTgpMDQ86RBnr6ePySSLk4g5OFDp757fBoc+Yhi9S+69MAUEkIB5IWNWJNZchMWq
/D8pnlHf0jzZfrHedQjsClGi5U+sJG1wszHejBoHd425vA1OQql5KhNry00rlWfbTP/TEI+VmseE
qtU5xIHnsrI4gytUY1RMIHjYl1+pZB4aYCADpSAAnvdgyZhmHM41QXskPrehtbZRBUh8X8rLbTYM
O54f9fmqvskZdo0IY5pF5B+VVvGuru1gLKhYDOxMWsxd4GaZ70NP5FX4QMGVocr/ssPNRjl6HMJC
1F176g8bnsA4aXv4gSrk82Z1Hh20irut3DvbZa9X1J9kMjrXTZMXQrC+aal7Yy3aw4vhr093+DmZ
sxF85r/awqhw5sFuaT3jmI9m7fw2Kql/IdjCYZ1gPRIyaIoJ0mq3rAeP6DFh0LDSVqO3F45srmdX
lePgQQgWkumXtK7+bOoVAMwJfgkwhOmT/w2imoyENbcI3cd3jZDYteyUpBZvk7TD8CyE720+jqYf
tK1UKFGAHqsPFkr3hHTmr0jLnMUA9Koy8aTWxux1KGfAA6Ro5vwc1+rM7srsaAEMLM+AFpEMXM0y
k/sXtXmSIZH+Urjj7sLvp3QLFhi3ZNIM2JvuUUQHzyzCi0+OZiX0KWxyX4CZfsP2jyUmz7mmanxj
SiNnOOBrozPR9mgCDP81sWNQHBXc8tJUfJxA4eWYVGovuIXZC/zv4ht40rItJAUCx3z+jDuDEwoD
tfBYjfGYrjxt+6IVT6HXcoiDaVMQl5nzI0t7HO5GjX6O+JpK5DVyWNGA75adDf+Y4vED13E54rZ4
SSmGMVE5TnEu8Q2S3b2zTgqYW8/rAYSjQQ42EGo4CqRoLK4NvAOoe//PtAItPSEoiecSACS3H0vt
uuBcRtW5tPBBzy7bQWVhLjuq2dE3btXWh7Y7LEBak8iB016IHIy60KoLLJ/fQw6Twdpj+MGHFNuK
2TB5Krg0NmIHVJKSH9221d5Zho1IShn8I+jzx22ypAFHbzDQJSXkDLHoEPsB+Z+x1RBG4//nIpRV
i6gYiaNhgehOItMHIozgWixHfEMQayInPMi4bato0eTFM1pabqA+HawPSGF42Ylype88hPEK6b5f
0/QlI0V6iuq/3GaXH5M+JVuLl84s8JunAbSqCNSKU1rIKHsE4Qv2j4ap0/OJyWVagN/6UTNjkVSp
fyQvK+ZGabUFrNyGl5zjhMwk6nF12YlMVGN/bZG3L4zxjhAbC3JYBeP5L6jYC1qrgB8wpoo9XJ/A
auv+40lcRP2qi+P0iNyP7cSI3THUNa49XXsy4swu2ADsJktL+gaa1I389dnUgkEMdwmdGvdTD71v
xPR+5taW24cLm8ffn/vmDgg+zieGxGyYjQgPiTlzbTZCa2kEp1an/l39sMemeXN1yH35jBGRJRUZ
BWqkb+dW80wmk/h2DBhXZkEGOZUTrzpi5u9IJYUhimOAXHgVLRz9/Qy5/BMVPCqCMQH9VrrbtFPP
FFddpUp89sNIj5R0srRx357kbDx2aeb69NRC9hvzxhGplZqJ5RtVa4gCPR4ZMsu3A1E57G54HV6k
ZOmFPIYoVcpO7k/gqjORflCg6XmJL+sguWdQ41c69eZoJ+OBvCSAbns9loaoCtD6ESggjv6G3r9X
7Eq5Q5Pr8rdlaMlEWnNbyViMNvV82ZKiaOkCiIMf4WcPP9t+YMwTIzhBVOw4Uy2HbuS0OV+60lyZ
POiVTGy6Mee+qsfktDpNA3H+AGZSByWOs8ett3m4xwNngQzU48/xl9chSVvsMMokwFM5dQpVBhvW
sZhUauYFviP9wwD6G8/APuBq7RhJmrFWxsryMx8WUACVt3vL+3/jbK3bd8+kYNPRiCR6OdvcqEV3
X+MW3ldhwfUNZLT4TOf5OwZZ5YF9f3joJndhkEb7E9rRGvC/kQG+Rs5y8cob5IwbAdjzuQpHGJfr
JoUtpq3/A2e6kQcLcLTV04TPs+J2iBlSj0ta5Ad5UxR+Ar3+jvP4rnmgJQkOWZJp415TftPu67ro
UHYGE/Lpcc5sQ4BGgPp9TOTWUlxxUdIi0kS3KLsTsMk5WyvX1je6vOphf8rJM7mhFtSOyIPbLbog
ZL2pCatXYdWw6lMnqxnXiHVXr4DWb8g0rYJOvnUxDNwUE9uakWnZYJy/dD/f/EphVejRMPQa0N24
sVPiS8VXNbZqTEObxPsNFm0gdD5IC+k9DHk80FFrToXdq/J+PykrRulNnVMf4XOofSOnBOTV17ta
aa9CoySQm54GmCeNMZXg6j5WJYT/JVFLY+FHYFmSycmXC1TxC3WM+c9N9/yyq+qnCBrdHFD7xTg+
6sNsLrFjauXJe0eUFM8OVNtqw88KG3sk34Ol+NOAXl9ueMNZPm278N5PbZkVzsyM+kNnH5DwoDBy
qDV6lg4tJ1JMQYl0he3A6mWz1ANqFelcOm8CxtgL7mvgfkvRuxbo+tf9qX9+vFfX9rvulrMRskbL
sZg42QCZdxF2Ni6+0N0qocKxbEpU9A786umRoyVeSFUfVCgmukxS/t6xPteSLBbI9hMtSvLD2xwU
BNPBSRWXw0oFCavCGfJeA/HlmJmlXsEdTZrChn0f7R4OM9v/j+gZUMuiQ2iMFk4iG4eBmpiIYeRe
xxG3eo4jO+s5pcZcY4PmM56x+gFLrAH99qHvA3IG62EngxNnJ0prHcohNBCRjEc1KofdTmFRCa4u
2zW1rlv3mOL7eGwEA2IzEnX9qKjTm0fxtDaEB/RMFB9R9OaA52ewxtcgxf29TPItFIICDqQnuzEW
SoBOYFXVmW4ZycBdEvoI2VxQT8L+Z5YvloZtVELdptLx1deqUXjbr16t/ZMRzrtuhqaurrDX08X7
nE2L6liiQLZIgX1Z8De+t0rxpcTXjgh+f63oanTlrqVCPam54Qnn/7WIoew3k8Qg5Pn9RyOoqBkj
O+lS3j276E/vj5jwDQfokOqFZBeAccdvbYCfUdTDwZoicNY5EZ8ZNXCivH2wwtzlE46mYtAhYTKX
rGC92Ojq6k5hveh4SvbJ9+23/hiLnzgvDMe7sQPY7M5q2B+dFmHxQ6Ymz7kCCS3Doopo/ECja5lL
BNtiPqXjZrytDFrR+Vmi7/vU1t1KZsGV/ANEcr0nKw6RW2MVwINAx9mBrtK8IJHj5r9G576IeNVe
SqJFX9ZhUOc4xgcRMgYOMMV9vhICBtscmZVT+3Iw3619RbLyvhRXQ6Dh12WWP4aIl7cKky0mYA0i
uT6KQu05XvOJkn2IeJILNGjmvEcimwtxsnOpL3SDSF1UEODaxxIBFk/Z7c2vs7dolCPLJOzNfqjP
XFF4YMK1bxKrqnZixkmCthOZr16YQ1qSF9H31UPrvMxdPRvMEyCAroxWITbEPM3HsDh1nXwgn23l
hbo7JVTWmjpei8Ao1HQEzlWaegP7tWlcFDytmDlFsmFltKz6NzAxzZP1ZyAWV4yRS9OgXkrp4WUz
7ThH08B8UrUhwtLS4E20NFLZDLyljwIPhirDz/zjg9nUlQepzNz9+xBiqusFVL3MVhLnN5gdNHRX
LhSSC+m1ejdAstD4kD85B5xCDEG3CSTGMI/CycJ00j3IRtH1DZCe8G4C+3s52Vp1lOd9vkAjsJt0
Rs5OkANUEyP240E+eMjs3h2rdFLKwYIR7SsmlgdvE34c7JOZqymK5VcaX4ARnOwcaEASNBtL6hWK
3tfGYSa4u12PYIZ5oIXOktfJZQU1qRpzHWW7gE6aGxB3gw6qv7AGB4QM71tU5UBUtwYMn3PeGJC0
0JEVWexZuLFAQWOJgy7AZlizKwVypc3oyk30LbBzNopOoU0ChyUAtTjdGx2c6ldNkKBs7sJXkxt5
uuCvd9FiWwxpa7yc9DvdDQrpjOzuU3IjiZrCom5+y46Rvp7TjK9f1raXMSsJ98+KGJC0U7CFdghc
sr4PwOEfRyRbZgvTJSPwSShviYBkX1831zE48O1o724xmcphAfRtW/RsFhFgWSJOTDDq9w2Q1HVZ
azaa+upJepobF7WoZJMpq6ZJiPRoVfNb0K2XhFqE+9m8tdiEdBfdrPs6eaJ7EH9pfEBfHNUjp9X0
TFIGxiEi8IECSLJONK1flLT9OdQiYa4w2tZQHEa0nh/KbWDOO06PYEzM8t1NQjLoO55f8Vb8M4pS
FzJMe0J4h7D7Mov2xLjkJKl/EmU3yNhK76CrrrZZgxLNAgJwb0HU8dj+amSX5wFfLqfpqRg4IhYO
mJT8SdAd2uyP1RXeilLRpvyn43zFmdKbSZ5Rz/4QdM9N+7RJLPiOaNct96vRV3GmM39Ty/MPQMKa
qKFfWR7c3QQIygdjFvX9PIbFbdsle5tITONwMZCHHLm30PvWO7Pd2lONEWCGTGIz+AlPhN0sLnif
6xsNrUnDipymCcCCvt1tvv8zWZ200kNNJmuGbrl67dxRv0umqDB5TF0eNOD3eCjyp0TKSG/AKFs0
CzX9yOFxHD6FgdruQgUS7VsOWGybcN85a95VE88IN0KcRblcOMFB0kAoxMhniPUnwJqSA2GuOwKD
lJo+kBm4/fgehMpYwEsYV8B6wCH46lImnZvr19s63qWFk6tWqxJUgy1hEdZQuXqJQf3NPLxQm9rn
RM7jcNnVhBqz4Hp6uwDecQcAwXu0dnsUzn0MZ0A5+fbQu4XLaiILYZgn0LM+BOKEN/OhW//lQ7UC
CUTgeuMZSmblr8MU7zjhpC2U1xWT6BKduuLU6B8CZxKyTm7wl4lcvCMuJfriFGDyCKL3jpzmieYj
U+14RiBuSqZPBQVcorRbMp+RsLyzXoD5ObXhMzViSOfoW/D+p9hTqsQfabgdPEYdHomYMyh8mJyJ
k7Di0L92WJsKQEJw/hpt69zGx30JHsjJ4oHYs+dAoWCGP2hSoBgYNJeqgfYnJGPvzcmSlEZL+7Jb
bsLjp1R3CdaLXtDi4BRcsE+nUsoGMqRcHBubTRtRc4s7chQ69ULJEqZhDVj7v9p+eEIErn6974ot
VntZcMt5CLFYhcjON7bNO0wtvl01AwaduY6jiRdRNJ68NeE9ZfAuPtvAFLU+glX5Z2qxUtWRElNV
x306OJoeGJlcfbC9et1cXFPD95DUMEoF56lP11t6Dlva3d5FtpC7Rlms7swuedbCt36/dW2fbaYD
WKyLz0ZB6JFMfcku7UuDr/cOv4Q/FhS8rTv7GoySE4kkLTYZpP4+cx/IF3HjtF061TI79Lt1EylA
AKWh1mnhpZf2r9sQA2G0kXPQWhuaGtufCcwS6EtiDgU1Aa+bqSIK5jOs+lucepGQXQw9BTqk8lPt
XxV4uDig5MpPaU1VFEPN4fYsfqhYW0niqoJl8w9gD4D+o/EwBpNi7v7NKUWXQBM/rhFzE+baUkd0
pSKpCiOptr1tUjl5MNGjEX5j+zX06weoFrRttFapQMK9bVsovnKYBkLWO9HoTOomzMBsXZD8QXS4
9k1rL4YMN0kSA54ZqnhjM/2nV2v797XEJYObosXXiyoJB0a6Xx7C994SiTBDo0E5AGLSzGVI/LQm
GrOucFkOAfi9gA84s9D9CeL1jlR4/lrPe4nYYIbjPgJXhTQ8XUkLDHDyAbinV8C/3leBP2Q4oe+L
TbYvYng9TJdY8tRihrSMvQHS6+DjSszci33T0GzJeNq3wa6MZNko1AHe1o4wMskt2MxhPgsHSEIq
Fq8usVO+TdaBHOixm4G9sOrQ2nafAGur52dWtooQau+CqXgpBmzNU5Hk9GcOzu8DQG4LB62grfCD
D43V2S35St52Ac5MytiIGztHSj/pXglbVPJrPUFGXrODv8FHbecOJYAX1sJxHuf053fX65/a3E2B
gUuB+RB9IQf8bcKuRW/Hu+dnjFyBx34XOcUFMMJvR35c/1LfG91xFdjWRMii0gDbQ2zaPrZIOMaP
KxvrWQBZ7BOZ4y85MhqPmfL7+0G6Wf9MLRpMJhTdUecP4Y/JlxiuOANfATL3Il2uDNh2zE83aYTR
ZPS4RPUgmWYRG/skVk0yjb4mZlYRSsWYviGzrWdQxYnqj2M3V6gEY5rJBIfckIfvL1iUsZgh38NR
G3WKjOZE9lDEzWSHtICt812IItSDmkxBdAbiJmvvV9cROZPp+h/JPKjwQjSz39yb6MGl8lnsxFdA
o7CphFhg81D5hsdv5PmwG0MCiJLde3+wrYzlmnYjrWEWlf0px8yKAW10yxfBD2oeCGc0HAAG6KOe
J+2jTXnXKUOtkj/aRt1Ou1Uql0rGF2hhJBkQTFL2EgHkLSBIywOfPuPhc9WeviY/n15/NF4EqvBM
cemo6aqy+bWdQHCVknCs8roIRG4MKiNbZSyEVBVouNUbS4sBpNCHTCy6s3R53r4SRiVRq/qaEEGH
wWrovUjYgFNPXNBuwB9/SKPG+vYFLq3jiYMmZpAdmxInnhHPlyXmeo5WnqWcN+5kdK07l0zWxABZ
L9sLO2y31rZPkiz/kduZYLKhFAJH+aDrDLDr6Gt4XbQumVBe4UmsTsLLfZq1WF4awCHssn+iwx2o
B51pSt801ICZqvq4O1CIsRlYNma0dwQrqi/JQ3rLv1yQK8tauEuFRY5Bcs2b/PVkYudUqZ7/vz7e
e1vE6Nu8H+cNZ35Uw6KcfV8alEI7IfTPWv6tM4d35Mk+rZ/UxUGUNOvtFPYVCVeRkFszxmxKIoQu
ksfZHVIlJKKPcT74q3Dj0+OOmo5VdcY6jEwkxfBmT2kfWRfsvRy3X8/6BZu55GYCmh8anBO4JVrv
QjaU+PZ+zxQI5pgG6gCe3QIhjY5jPYKoUMlRWdYo48BFTCYB//98eWUiXedqBIjxHBj/0YJd+lIn
3LtkADh+3+Ow6uEP52CIBaUl3MS+mN/4+D2m/OC9txwGRroDPKPsmTPe6ET8rPdDTHJXhEcstjPE
qROxgPtSCWaV/55UIzyX96aICJ6Xt5l4NrPxMRues4E8seT7bdqTZlNzwAvQWSNeReJjFcteSGUh
YCgCEGF/WROR00SiRhWJBF9EigE28qCicsUaXWJrdi2OAZRCWCYO+qJ66woxrpUHFYakhogYUJt4
88XnasiOLWwEB7u+IISBE1/cMKWRt9S2S1LIF+N4TgTFEXmoHdXO8/qVLYuy0bATmQxIDb2RxSyh
h13N0+at24/pmErJwt/35U+8HkFWiOy0cS3YB8rTemncQalO5jyLTMQW5UfJDEfY6wa3CPKekW8H
axJJz7vifEFD6EumnC0YrBzGLCMq7Tjsk+6Ty4O1T/2+9+Fu4XGRuaD9a8HB/iHuqULJw4rlx5u4
KxrO6mACfVx1TZaZfll/jktyu32rHXkBlVM0iV66wDB76FZF51/Kf9xXODDgdiTyCLFoLHac+cTP
CiHnFj5k6WIU7kEcN51GoX8/7WAFmNI6AtJF9EES/86Dl2H6KnC6rsI268BjB4jDhFa7bo5Lo3ie
Jn+E4BAlctgAK6JKP5w1XWoVGTMn7uwM93ukqpPrQYaDajKq3QcFzDxPzp54lRrKRNHbmx095BFo
you+rLYVpjZhUrfVugXnQZH0B15ZOZ0Yaw0wPzYnfpHxeXABRvRfBglqLzlbKIiLsYPnfQ2EeWxJ
jZ5AkL0MES691Ev1ZLA04Bd33sh43hqxIsvcrDfZVC8LOiu+babBz2hm4gtaqjAN25e6NDNq9k6g
mqxLGugKriv+/q0/YIiXF4QmabX/nKA1W82l/YIsdWMMgtvfCthSmQgcaCs8Z2DwnkRGFc78lMGD
RZIsTzxZ39fbudZ6uv7IQXMjr/ZXUV9A0dHUe8Nx10/4XFfkqHncHd1imMhdFB+564Z7ugompk3R
I5p9SIBJKIIR5Xq4sqm1PqOCDBoRklWI5drlXX4uEQZr+WYy5nYIQiClh5Ib6uGOciFl4aMkyFoB
tEKPOHZmYLf++Z+vKL6oDriXGq100eTpaL3VbCDkoni6uUCJQH1muKvKv0guPHb9/tMo6AAqz0Zo
FDOOgGqEgMjs0INsgPo7etgRy+NFhDz98qwXm3bhoixjkJXV1F9kRrfcWYOjyjD4HpgvZ/LNeik1
0RZ67B20xOvYHBpk/EL8LXdRjvudgwDPm+sM87qz5ClijYBHZ/wkqkP83TxaH4frHbd7THpjbCZC
AaHtdVBn5C+MQ9m0NZ9SCH/hon1xSj/sW7VEEpvll1tXMRFIZUNKGWIGnr0dxVb05CZQS1wzOF8g
9rza1nN3tSHhvXSZjFWslKhifUAEFhwX9JjgYHKfx8EXpd0oFG2s2QgwSqPi5aUlRRd+urHyvVTO
JOjI6kvsuAbniH09Y8N1x8SofjKKI20Q+8xNSlrCCZUbQH23DyveMl1p6Tp1WnGHQGojBEKaX36O
JJ5W1IjJOJ4UmTGgSGJBI3XYY8HtkAAAR5JZoDPahgWdRUxHlUWcc1lMqS6KeL75tftCYCsEnk9B
vaBlpC0G50VI9sMQ5xGyTEaltOO1GIM/PFFBm7fob6OqwLIMDppj+pZG+1lzREpXKGI8jlKj3bot
3KVsMlE5OjmU+6aYwCzeVpjv6v3LztizjLd8DrHUAsBYT4LIlbjAGKZXls6ZtVElzLZQleOPiaqZ
X7ju1zqyhq/I7LxUDQNkEmOYkbwP9aoSZfqA9mKHuGVX2riULicg7wvVT8oXrqQevKrZLmIesoMg
N7MW7Li0wbCWvehFVrd5OAkbQVJsy5C0zRVKqrlW+rw2wkcBjvMTOGc2o+A2jL4+oMAU6veMMxGv
/MLMkgO9dvzlTBXeyWPImTFaC+OKYHv92QNwlxsjP42ozH8VCGr7ko/1qH7USU6R/+l6VLZPn9Jd
USdbUAV74FYYKdJgErsKIPoGyJVh/SWbtP17XKk9O3hjzaEEwhRS5xYi4AeIYeEgIxl7OoXf4Vli
4vVxCiYQLJE6bvRKABChj3Y/COknrChk3Heu1gEAcmES2ftDDfM7ZMVPLQx0XxqoIkP6UgxAxr4G
ociVCRsa3NZjrw8TD2zxz6PLbx1184kZgahBjYzQ7WgNr0NeKKTMn52Xj7IhPuWRUy+CsRB/Du3h
7/z8I9vuF8AmTxl1dYqCJhkZvB/BqAChNfNiuaI2eaBRhBUvcVijWNRDluaovcMq6Kp1/BY2VBPy
6QA4U+kT38+Bu0kBVe3Vs8dtRTPuQKz7Hm6tJTneuAswfwL4B7xmd3/1/N/GINKGsmRg2UL/a2J2
eTmP1kA+ACy9GYHaqD+JuT6JV7eA8uN9+4YI/c5nCUz1ZEE0iApJsru6XRrhg9uERLEq2CEXLBRe
gWvmE7CINyngv+1PC8V45nngLpHngoknCCArAe1JyYtxi2IDkVsRiFxDDgT5IhuCmB4PPrcMa0ay
YoiqJ8xrv1OWCw3m2RHSP1Z76QyDU/bJb03HQHYBYcM7qO68jG23iYu1i+uWgCZayZXmN55Aww2m
3oD4Mse6D5BwQBV045E9XLBUI2H0BlmUvAL51iFGEmfg+XXOdwKd3o8xkpDt1trSfNvRc7rknntr
ngZIaPJ871T21vYod59SI4EjJCHw5sXqLXAVWdxQI9Zt64EvJRI5gXHlFOLAEo07da1q+TxUleqQ
A3wUVrgx7lj8lcxu8HlfnLJlIlYh3IxJeRRpEu3sBmicRKc9pmswsgdC0z7MNKNEkDIDmd5W8vEo
TELK2SXdQec8juFDn12m7p+fS6UE/19GhWzVAQORm6UaKse4lavSPPyXFyE08egzCkLUKvv+Sg4A
KNnxiI86fTXsP/vrwDfjwSjAWvNgzU51mkl4V7q/ZqwaGKN1bjBsQ9WAHFV1VEjFbljNXCdA93eK
4b43PgzGOBQ1yUDrHcyLi77g5Q0OQopQ4HEdLRXJIJnez+e1yDmhs3G8EUJQzqDp5IcST4ykUm1U
2qEGVwxP3xwHFbUtYUiTtq28Fx7Zr+WnMWXBbegxMWsHU2B2x3/BMnVXklQ7cr9ICqJe6UjN0lFV
oHudGtfD1TbIzaQRWwCufkM+38dIRF39MsA8yUGBaSc4HM7ZXBtAq6SwDxMJLFLNC4h9oZeeIQiR
70Tkp0izOK1NwkVWar/FtMHiSrl5ozkaDjA3mM1QImmY6qWXCBn68lRY2T1qRN4GbwJ17ijqi+Qx
TUp9XR/KEnNXuf/A/WeRxVzjSn1W6ymyPOUXc8SwPgu2HVsXgtlEsx/cTstEehS4lybd4tB7Hqk3
FDpQ8MXMNT9XReHPr+XwB6EW9ng4VRpNOOsoh6ZH84TCpA4tbnQrRRNyQzd90IFI0Cl0ojv8ZbI0
s1ty5Bwnqtqkpz3DmWVyjVxeXWYLwKbJ3T8ljzrPfqp+WQJ0qTVXR+zkae8t2mNaH084IF/GFbXI
Sb4PjoDhfdlttVhvnGbxReaC8pAgOjX6GzphDzKZOmph678JSV/mo+q4rePgns2xDTAcGZ5jv9Am
OG1zKPMALAfwYG/rj8/XHiSN1Ukym2lQ/HczhhQD+Un0K7WtsjS6R0ECO7ufDRRpRRmgX/rTN53s
/FOpefMRk4PMGGMFZfR2g/oJNyzOlAEL8CljR3HJyf0WHLCwAtC71cKaTC0FKC8vwWwrFHZh/Uwx
GvGBnFknydo00UVcHaLS7T3+Lj9OguY5qNrIQVhWOjYaFX64ATd7jU1tc9FSA1ujzBnztHsFNmLg
Q5MjzWV1xnrqGA8bmiYEolZzGfq6csfEoPVnrqGPGwSK3LuhuG7V+SnK1FlsQ3Sgwz2JodupI0T8
nFyNs2Rfd9ZLHnEF0E1Z+1TWhpARRWbwuhi2alOBwS+sTfuBtaqHyMefn3Nw+8fACzwYNYM+rPTF
kgNefPg9MfSqFnBzopUNJCju1XRv+8V3sqdddSfqd6g2qJPIfbrX1XUFSL+DywPA+41eJokvceVc
FO3vY7Rp7d2uF5I1DgnM3ICKFjMuSzyPVsd3PHaNPdq2sGKVVMMj8/i+M4nMoTpyBSrfxffY6ejS
/0mm5UCiQiNJrDEMYKU7xp8n/GRThJtvfQHbaXCZOV6XbqOolHaWhHezHQpUE3XObpX8ZoGL81nC
0RTMJOC+NU4dOzC/FEV9XU305CSFvSqNZFIjU9HOFjrj0AQm/QFSUhjppc4d4JEQKI2/96Zkk1mV
qoIQO9oOBqNgvdIhHRELMASpCPoNGHbJuZGTzsIEjb6qM8T2rVz/OnnxRYAgZdhOx+EfbLkjafIb
JpZSNPcOa+o0KRILhTXobnxiDl0Ia+VZTW11ShABzyD7Ploq2v7a/gZdzN/rc/7AEE9WUe6XfYKI
rq6os62Jhn3eTfAcqQGHJqyD277wkXELpEIZx22EVaoRc3Dc9+zufn49fe9qjgA5SK4yqFnZluOF
pY99LCf04+h6s8FC0A96Y3QwGxj+NRecwVfhBTO5Wg4h9K5WAkLvcMRPrS2WmC1klyscTToPtmRa
g0Z7i/DqsExoXqBN28A9QoIA77Gy4/peyXQS6UZLetvDTMPawTv6LYmZuhnBvrqWTZA3neWJBz8M
i5kRWxw6rRpik9KRAupdv2S+KDIrjNVJ9f0aWTTM3X1TPNKkUWtBZQzFGfw3JoP2aZM+VhBxJEWV
Lh9Vom28jiM58ULaYeWfGjRWSFQlcqQ/ydVBmQs9PZXDVTgr0Z9tdlDIFMq0inKSNU+TOK6PhZsq
kbsx7RWk6vQmQsKxK9qmFVpSnTl75MYVTZ/HODLnSkljP1fIVxafqBC5HcMZ/1WycpAfkmuRTFg3
Vo0BQvWg0ycxl1p6XFoVCp04DmTUQTF5PsRWq19TjAIDrXxffxMq0uHK9557fl9uB5LDrnGKYI62
4XeJaeEAxpCLKJiJBCxmNlpGZl36G8m8wm54OBNe6DmQ9EOF6A7Hx+1tiX+1L+ZuzeCtBoQig4ti
ErYf3w7zKHJa3WMcomk/Z9nTlmAuKLoW6A/enDHzF1b6EeSMzc7tL4cyvRiMxX6dgcKL33/898rW
mKKQ0qkHUIEu/38UTeAmZXexqm9bpvLtxSSLs6S9xLT6ombHVI13bfkz4Sg7BFV4UMPM2dWxw0ty
J5VLG1LYCzZII55x3/tPG6DkTN+5NVNH1nNXWYdFTVVgLqbuVkleo9pymO+sijkcas5uy7gPCXbf
vCBxz5fK6E2EBBaa/b9qbS637vl/kWTtWgqv9jRbdxFadSDtGklBDLc62Nhqk7C9rvOQ+htUBsta
zROTc3KPOQdQjuUk2rjW5Ic5OfYz+3abHKzEfmxBqec7ff2P+r9Q33IvFYa/BjwUgIXHQPoDQMT9
y8+pupNorqslUBf6RqQ1B1kFFvWS2woTTddjtMlDgz2LKo3WDRy1OBQl0UcT90+ALg3OZnh95YR/
uBq7+jtFxxrxydKCHK0txAbj5/j20odw+tjUNpiX9ZvhL13FMDuf6j9jaIa6sbTx1+45QGhTQyCt
2f9vs+tbNZEG+oxiwKbVEJCfWJR8nKofeGHGorohWdVMj+uaVCu1lK+WanjRS8I3o7mmyrYpjc5Q
RHPqlL0mq5aIVGGQiW3oe0Hpi+Pqnl8jFZ+1CJBeklpOc6ST2R4d+BoQo8rXnk5btiIIh3xGHyZc
QdLKlPfUgKw9wMVTXufgkuNdRtDE990QA3K90GEBGMYLrT1qOgNjWuw6LxZtwEwk6cDoSXkJhKrE
ifwt3WXKiBYDIm4GhxiMJqDQwBpTSMQgl03usSMFOt46+/1ihiP5rdJooOHWSH1xGs0bETD7IfYq
lSEdI7EHCHM8ofLmRDOZ8uN/ws1kjbCxtMW//3aFERqdk2jayUw79HcpOTh1cyHGzIsx8fO7BR7N
p6ryDFkmeGAGMgPge/jMGVZMPjZ+XuGEWHC3hyKFWS57ljMDu2TR1pDSgA49/43VX5bZ4UUywtZ6
+sgp2ajGLdarYvmlwG6JS7QfCKTE9xosfgj7YNoZsHXrRnOCmpyLkR4G/8nEf4GhUt64BP7qSXSC
lIwrIBZeG+XbAzAJpgiZYkyxODriMB9/vRh1XoWPeQQeHwQqVlgrPYTdlI3cG3pYjp/f3nDsJAwG
0wtYjj7/VSQ/hH/hpSzrgaS2OaxlqVC1LXF3E6P/+Hc4gnWF0wC1Q3sqUevMuv3qiVRCY5Hch/4+
7B1YB5PPduGwytQirKh/y0ijDQudSeaFEMvqdO3ZOaXmXhRqcVxWpLYjDYHKvPhp/9cifYDVAcNy
cyyKdYINDm/WzRJ6rGtnz5bdA+UNqXE5zVcigpSJR0HPndC1vdpOXR9zTQjfMRYKFwG9YC+WURCg
5+gwrWphOnELG3d21QzhDTPWDus7FSoAz3BCYMJCEZgaNPgwCpm8l9c1RQcJgKQOd1TFNFlDigXZ
zlO+0hYjwTn1y2jN0z5eM00AK/dRgGQVJwzd3iZdrV5/Z8PPk0xnfMRj6Ztd2mGOOb3PmlNs29cm
+eblHjK2s/55Y4HkU4CnxwEF499JqU6ySKyV304rvv7Rrk4IyYinamyjtS43tqYCjPZyw9aCb3fH
kkyVpTtGphWMQxu6W1Esoj4fD9YHQzVpcMCdZeNFL+3fl2uspy5QFOi6YhL+FWJFuq76/GbxJ5+t
1QoiJyTquw7kamUpy5kaNGf2UfDjBm5LTTLmWaxVS8+Nqiv94jxRULm9MSrHFcRTBkmA1oIr0GGU
BOGafVWtGTBp68lE8LOTxtuoT2Ne1xbNQyBCa+nTqUZwcexthLae4Nm09bMEfgoLVIB9frzgRapM
NlEITZ8BQU2GJlEf80WhaKzgDSasftRi/f9pesZ12cS5UhDQnr9xQN+uYTikYfsHVAzZmxBGwTrC
ltYtHs3lTUz9TnZtJaVA9+vpEtCKEHInP1qkx7x49OjNLIGhwa0VbN4fsf4ut5TQL3gVnS83c8bC
czuZ7b2qcXtw4Y90iQmUKkFhJoWLjsTRp1jfZHgW+bWnsbxOVTqWDNU+FR2m1b/m7CgqmxSs8nIu
LHmK/8mdt/d7ur3VURs1jel1N7x/AWmLlbC2g+v8mWAjyVcXtTI8LseJgj5qQR1swaZafltO2wcH
ZDvPv0GWBHzyoA5uWcvR9RODNWIvH6yCadpTJvR3MK1DDeZeT0wa0pBSaXZt3++RiK1tXWG2+4CQ
dYbV5DV5/cRSZzrUIN3iJv93VChfLTV5aToNkYWK+KivtNCRPua4m29ax81XkNlBLF3cho44bjPd
14r6NQG8ltzRNpncoIlOmCYFAre89D+ocZxt+f6WVxhEzfGZoNx3exQm30cliI5L7A/RM9d6Xiq7
auykHEoUv9xLY3rJFnBIx5wjTB39nv2LjsjNNqoWHfes1SKBJjBVEonfzmFEAP0xmqayMjP89vL4
ZCDT0VjjEHcVpSqtpNp7MXz48Khnb9tZsIFEbbQmpvyH974LnNCvb2aqcM2WzK4ZFfdMqcPbjvVs
mY6++kM8DcEqn4TcIxr2dwkHPzunTU56mRlEydrNqesUmxWIc8YfJG+0E/w54KIN2TQ80UXvhCZp
JgRnGG3W0lTJZx9iq39iFgE4kkPN4Y5XkcL/rtAeQFKSO0iSQZW8iKSGOPA9Fpy/aM7BKx/8IrVM
hq+kRT5B7rIY8EX0C/kLXr4Qs6Lz4hiLqOn6kWxMzhAub46mo2eLQ3y6R1qiCFgrkrbA6fELHyp4
s547FSXlCCza55aR4ZcFHyUKdyoNZa5WPeBriYgFXxCQkqc3Ny3Ip1S/2eW69xUZ0j0LCdwHRjF7
pCXLGp1k+KK3ymST2YT2AShLUQ2F9XqCkWKcLbrgtZIBHWKfLFjyicNFzfuXevoRXZKUhuCR6DbN
B1VPQa3PxiAsvHw6pFzqA2zjSPw16ClguIt6SawpYS+rxatJUp3xYewBGjCqUi8snw16E53Ebhs9
0vADOmzXEivlFWDRoJreUfb2tqQnDV+ZfXDDhYxkocIIKo11SYttAv2XIkoaFGEY3UpKEBwnFlif
Qd687+l9vt7N3LwAexgMy0B9/91zmlyRjO+fi5OPriN/LDQ7EHZ/qg2mMcLV1yVQDyWC8/VpwULo
jMTJQ6BKSS5p8JKTKNauL1Viedw5S8ysFrMJzM9sdI59IC2NJBO3PpSWRHjSsrj0RMp5tTYqo4CP
+bJIKaYW3kznxbSYCLRcbIpc/Ldw17e5ahf0LjjYVB0WK28ncPUItGq7wugP1TUsqJw+LzW87oGO
e5JrD0mf6Dn5GYBAp9jQ2Ud4hO3SgLDvgaXDkmyTLGpDm8k74qHFiVvg6AcKUKTqN5Ni91xXYnhh
2wPr76+sBKQ9FVKywquq6ms3mVVsGABOcqndsnmu0LgfPQWvGdzKv8/V+dUeIbmAtmK//6LB6HGP
ZnEqEUtJvmPBJ2QQO+LOTjjzZXUU6b3b4/gXl2nSVxz8eRAyRvOtn/GqE4XqqtXiDMTOi21rEW7t
/lUob7a88SnZYqSY0J+xP1ZemNG8X77b+VRl9ofvfX3glyNYhmsms1zKWSBn1m2RSSNbwNXtPK3b
v0oZCAT25MH/qdAZH1dROaNWJ7lAXZJfaangUgTCIyHmd1+ccM+qTzzNz70b0c4lq8fFO7rSqiFc
ZD6AR93jbegOrpmh8pCM7obGoYUc3CS/0BML8Msl42QaD+VG31pq+RGr+OZzMCKGsjLu0jU99eUV
u98LLO1/yQ90vL2cHZffwGI6SuLK0BZILIrkCbkymQ+QjFK2T5n3FwogvMbyzK3L1omjmzGNEnuL
yhEfYif/A/Npe7eyjKXx01wLnVVZLgOrpRfLg08ceC81PcsZtnx8LaDT60o2WR8+GH1AbI0lfGCz
ofiYg0HJVfFHOQgow9du3bqsUpD0oFAwGvDLL3e4kg4mIzrnsgT0oH4Rs/pMbwARDoqNGaSBGa+j
3uxHwtqwkJgaeZOSglY6xQ2MYYluJqesLyZAt066F410VXIbmMaws2nTeP6gYmeoIMWo/B8jqBOf
h1VrzUq1djlJeTXBui15UOnjYh2g5B9g71QVVNc6Hk1C0DULjLa5zCw6g/qIzgNFwD17nNNTPj4H
lyzzQy8hXqOiQ7DuIGBHDgjLtQnEAWGK85Rha5IAA3jUEktbdb+tdPbqRCPDiBv/DyQjD1EPle5S
zMNo3s/4g0pEgtcltJHJN+mMnHxm8sPwzp4aZzk/U/1zmaLoPbmYmuwcih6Qs4XWGNfEuhgufdGs
SFw3M/aQRNfsVNad0BjghhRI1y4I5Mq0ZpSCmKot7Zie0/p75MZDoydGXJ2G54q3kHTdmzenVrRD
BbO/pg1Nb8h342o4ORFUJiuZu/2RoSkC8ytXo5gEfnasBZCUBssVhMgjg0OSiOhjQcFmOSsVabvf
+5zc3UikiUzoTADlmm8624PJfOlLNg5C/kvn1mWy3mpiRNYSLurtoLFAykzO9XVmi90EYTfZ7Hc6
7CEfkOvX+frCpw9Vw2/A63IUi9PrAm3mTlnoxqZsYfOgEGu75BJl5TCKCQVOIifDolj/e6CGJwnI
8ZZT56Onn9c5LdCzQckXhX/tYPxQwSALlaWgyRvzlLVpE3dBDTNY/5jkUaWUx2bLpSa52GeI6wWa
33M40Epz6YU96BO/R9OxBjEPfnsDtcMeZeVHNcHu2xtwH+AjmE3vnqksMiAIpS3QWmg53F2GbStZ
vlOjK1VhywKLjyxqoqLkuL4tsscLq1cWKeA27lGspU5Gpp7wsojfynY08l6c3m3unqMEP5KvGOCt
nofr/iMb5ZQ3h3R8Qvb8EuwOxLcEMnZxKGSEUMw+J7LHhZ3nqLIdJ3qvXwpjWYpnzybk+KI8Ylub
lSbBYRdi44eoK1C6Tgd74FvoBMqvkE2jfTSiHLJi5nOOYHk3tGdZbXycH133UnT4GZJ7DnyjQZpT
AbUIWd7CYCcoe0f1wEH/ln3u1zfQPbWJYKFL7Dc+wd+KpY7JklhuElysde3pKSVMCBybk0rw0gtD
uki8y67vItWkPZ0vkBHh1KGuZwstSPAqtjRIUx5ORZhe+UodCJiM6GBBMrVveBusdY0ooiBIXL9U
xxLcfH3CZqR/7XAeKodmDwsw/OcJzVD6Q+UPuDWsxNB5FCnq5T/Ns2/i7QNyu0kf1ZQLVPcoc/Dg
hxVtX0iQ0cS+cDJXK+tVi+AMmP6P6LJ2cRr5a5gHzLJ2ykNRLNA5NtdcfBN93ApcdVnBEZMVTp+i
6zm7HUOAO5svQodH2XT+KE1xWkjQ6W2/9h8LkPY9XfMlb/s69lC68Yjs8e8PDHUpuH2uxH5bd6Em
E0+Q0WtD7B91ed7iLTB3gH6+6lfXFu8jiculGk60z5qHFh/EEDWRrBEOblQMFUtZZ/4CmEdtXLXS
FuHg35DYRU8qqiZKNRO8oEPg2MVCi0AzRWBzTomXRLIDzPX/ctxfUcxbIslHHxPPhz92c2YiivkX
29hy5mWGHkzGcrMewp3sfuw6WtYq4shKdRqmflIYR8p06UjqYgvQdjBkwl05wYXS2jj9oqSAgx6a
AzScsdvhJPvgKS/tfUAXftUaOAKyfeRkGpJAyrlp2sB3HIX5exPm/ksvsUIleu52uLp1QYtNXNvG
mLMObmFjkLDsw/jUA3H+ZOebuurPI0dFBcNSsjpcR5dofgwxcNukIBTPzjWmkIhlkWz6Xdlsbfuz
4NvDdqhrrO57pjZOLIliWoH5syOSGE9MM145BMlU9AGWVTPbYxt5Yn1lhNKDjpf1hLuXwj7jyoVO
d8piaojTaIvufcM3dW1qGfCqwHAsxhYK0qwuOXY9QDBNwdWRfiNpfVJikzuYZjiGAxFfLuo2OGBC
MRflfcKHeubHHU6nid/N2wpMDJP1L47LGKL+GNapBSUTcR/qS9iebIL/OqaOc1Ny7em9rjK0tasH
krVWkdjSA2Ee+RKkTvb1FebP/vNUd4jsdF2NMsCmCvl4gB3mihLH6sNqCvmu+E+e0nAPS26xhXyJ
xJYNpxvdwjraQD0uLzhbdX0X9t6/Gj6BCbOUanwtH97QjimHs5sqBhBRvRYJt+SWjD4FSe3NlqqZ
miQagmMXBJDT5kAQnJLqyB20DoFa07pExv3QwUlL6FbG4GPlzScNDKbKZbHQT9nsaXQDRdiDDcv1
HwTtYEC3daDNpzD0W93PgHEilUAY2DKK8s07mg32YyOOvock4sUge3LjQSYEOEnRqUDbsiiLZGCd
Z3Q+7Kf96SMLeakx69X1IZeYVvnwjmOXk0aAv/Dmu4P7NRzMiEYa1JgwuKnCJNLwtF2wd2gr7l0Z
oFR70sW2MJnDA87YbN5EeAGy3btlskym1+Zv28DM5HgTdX9oEzojxM2kq5Sndlc7gUlsaX0et7jA
8jVFFfwEZXd+pBx6hnVSKeNswTXoNHz1prjCreH1gihOLTH8j7NXTOFD1AESnIY5p6ezoROO+opw
LdR+vBPvs2eAH10gIxs1KC7M2OzA4sy4VB08PY/kQCcnC2U1p5zXDkGNAlRaihyW6lvAZOMKSmb6
9onCIpdvnPMRvVSofAuuabYHkZ9HIP6LOytfCXqQvdTGTrZAkTL65MOcJ7ksKXtRpRr6CIhr2aLu
sjVoWSDrlsQ2Jrs0sc96db9hAo0KQOam0mY4vPeJhv32HNgZlaurZtI/TmPfCM4rgFJOy5/HPUP8
/yDpq7+HlB9lUbDjYC18ZQXVi7sg6A25eDQM0Ha1dyWRN23BPF5M3NXsC41CPBZsI6CCIAOP4CpG
BoyCx62wM9UxfCJQzTG5AHB/Wg8FbRZKTH2WhI0jplh7GtMFehDlYYM6sFyox28v2eBmd/vQ/w1P
bX0HzWjWS7m5SEXhT0l9Z3SQhkmclFvXVAwpMh9wnL0NT250MhmI/bIPqOCSSW/5B7CNjIQtcibr
CFyCA3bYXVzYH5vrTuQx2WNYJw32K0qpIfMRVon2xZi/+Z/X95SGG/tIm2Yxy+mL746hUuZDbdc7
q1RdeihaBIOHLzIY5mG6Bn/fh9aKObRg8oeh507EJuZIY5C7cW3QjgHFe1CVPjP1lwHAwF/w5DWC
lIqyyxxxc2e5OtICMUpsHfcUCKxyzsjDrkJ1Y7JB1ShNSbUxq0qSwaZkB6FOf4kDuNMAw/DrpU20
o/OneKKsciiBtydrz0k/rUyzn4iwmCULkFp+fEz+v8UW24Z92GiK2OeS5D+nXUbSaMO3Yz+g0kLQ
Kh3dbsxRk9vzIy3M1HlhQR2LAA/fhxXptDYE58XOsNpWXN/hcTv+RpFhyw2/3DDzyhpIlqvh8cUJ
IbdKc6O0rigP8lP/VWhUgVlqqIUpmayrsW6mJhWbIn5Z+VqJD6iIgVYggCEGooFuiIQdYWASuDSt
d+7zoyNW5/nZy5K2Rd72H0hrdohek5l1+ysOpsP67dsanswSEfovOMERmgGUjx2fBfKZFMrX2MaQ
DDM5vBdm2MAAnTiuzZsAC3T2SozsjQZC9EBruz6r02p/O7oB3v1IxKE/+H+hRiym5oF9M5blsyTM
0ieyx4/D7Fb1pi/v2bTkZSBBgEJeD+ZkgO7aWayi9zemVdmgzs6145DQdNn1HLPW085lxUOTd+Pu
6XVXj1mEAprd4PTVpndLmFReSRcLDXF5qhLfOZnib3gFKWJI92NM68bqeW0slMjSRRXu2FQTWOkT
GQf4bcMDk6Nh8YiepDI7pp2aQCG2CYSY8Ej9r8GWNPQBxgKe4AuJKTG9Eh+fE0p/KQnHq0H1ZPB5
83F/OMOIsaejYXq2LOOJKUaSBMrB/GcLqgBnwWqfp4wDklUHOAk03HZxl1pCJZRHgDF3YDgSrDbA
5WVk/6giC9/s37N4yqaai//lYDqJB6G6ho6vQRJ9I+3N7JruhpEqNaoYF0ChI/mB2makBrUHtiPK
nnfPkD0WEwo5Z8luizNsKeLeL9s3rxilg2W74Ht46gU4u0O2YCzgIx8OmkWa1YACdOZzUNzFaiHi
3f3oz4g7w/Y8ay6cU+9UeWyP5h+e6HVAo2KNbOGLQ8QFnUETBG2kBjsK18yTGbkABdWTOQI/5o5P
Nz1xtcZAJKbjmhWm9UtQLUVxFbeuqVwEVRVtKYCo+0pqnaVdFof0wKtG5J5IIcG8bIlayvqTR8pB
JGpTY8MefP2UnVmJbRx7Gv3u1k88w25ldYNfukjnOaFxAI03ICXPC+nwMTrPtsYKCA1VumieO0Li
KpUNmem8Nf6vMNUm1gBqzsGuqVDe7AovIK4Z88ItbsTVeB6EtvxAEj0AOQ5Taz99XN+N/jT0FzUj
M9LgDDG772kYQ4HUOC5ZyzXEC6XM3FLpgiRIHr2knGrhR6IBmxUAOi3gKFVuPahAOdxjIrjIIgXK
R9jakYJAoZu1ie+s2maJ4H40r3HxCpv2+dtoy2sUKXJv88n8Wjds7jFX2tLmfE76xkUXZiKtEGii
LVsMoyJWfN7VirC/HZnk0Xgu5YBjWLKo32XBmEseniT8/PzyFVpkG0EaMdB0OdxV8EgZdJmziZVU
FgVYZT8qpMKew/86SA/rJuQdfbOZ3NJyVY3K+gnityPnRu5gaHbHje/U2MN6TEoyz0iPHY1Q3QML
DidxKRSx+aP5BPxkLHa83lSFwh+sj9V8RwNzawLM9jar2RM9EUHAxOIsN3HeJMVnCOcin9lMTUIP
dsiYQczZLU/vMnC0vXrsTCAVVsaKFnwgMtZj9tPu3ME9AJu91+8kST4e9WBuoGALIEOWyTb4n99g
YMHeslhshYmvvayl/O+igSmGU3UK/o1ClaMNJv3vp/Ifn0RB+OorIBrllorQ+cqY/odpyOCE0uZ1
1wJ9vo/XNYzGEoCemsk5nNrz1+mKIEuma//B10ge9wshHxKpqDle7/HV8CGm8nE0EoiIYdgicNGK
X9Tfbhy9aMc2Fv4evrXt4vZ1A6e6RIE6Y6NKjak/tOQOXn6/kMLBo9t57MqPS/jwD+uJ8qlgmogs
kLpcvrpUYk3p3jyZgf/EE/U4e6wKoCMHdQUzHdMPcF2kDcXmie1mWtZK5CKXXPPl6/yCvQN1XhfI
8W8QVhuIqc6ANkV6xnnVsdpEYboNQvuJl0s1EHgpTYrlqgq8lkauBuwy0LIROsHaexaGmOTn9PQ1
fqavgp8jjU7S9mJTj4Oyp/Gvku3kZxSOXEEFuf36Cslqxa33i04bKuYn9DI6tDbZQ6CYZbbslhFb
7liixP50VS0GRBVyDoUb4MLkwlF0tLSz3du/0x5Qkokng/OlHLuTZzmmqDGbtlfvghxVQ1eiQ8TV
iGwFFada0iADRSib92MzZ2wDqR8qplc3JAS4xXUEh8H7RqGc0t8SUuD8qIvTZ90raDvvEFJYN0tL
oOOnbMioN+hYp9LQdWv1rm9LGOUfsy8RJ9cU2qeJXVIsvtzprwsQgI4IgqSgSIG3KRo6vWs9fOTg
zsJdVxkOAXWSb7zLrRJD8kge0QFV0vGcVE1X1oeltw7AbkhA5UaRlBQrgmdQPlMfnKnO0GUeBXdH
EvI/AS0BbuseWSffy78k+bBoC3Az7W6FXFYNjuNThiaP9LVZ77+C3w1zthnXc54wkjfHYAkt2NnI
fBl/dK84zC4L4GUUXWS8NkvY5BhLEioQdlSBj7Mlj9rfj2AkT79+/J17fI4M5qGsutiWRpr7FLf3
+pIcZmZZRkjqJC0sfSHLyxf+fVzfMlN0s9Pd957kyx7hA+QiFiUxIoDP6bZVw334eRUzvycHxttJ
EcL1nl1BZWR0Qy2CojQqm8OZ5K8QrvLkHLdYgtOmBFkbyez9cME0y8yKTXvuCoQJzQAzYMv/Svd2
o9uutHWjl8biIkrsa4p0/yub82xpKV8PpSW22ak9GZ2CmPzRLH9T0A7ct5d9T3AaaGORuVytR8DU
OGYI/6mjUuc1KosZodUqWbU6Omt+DmRuRKnHFta633lkhi9TPZWOaxxmEn1tX7LITEh3PAaYtQzz
iqRb9pI7gel+GhR5zGuE9bm5hCZKFNVgFvuEgvOS9JXgiF5UCVA4JbN2AVwqe+9TP2l944ZYCTKN
dZvuyjvY80pCM6I0u62Cfw1u0JGkinErPBC1r7TBux+KGgegEgEZpM9b5NateLCake458ZEQ6WGM
iYT7trSsk+hTn+HzJt0ZWeIBA5KtyIS7Nqi0SZGl/o1kKrBU8PzHy1Dg3ktHOFS4mvqq7nVhcVBl
/ECxuecVUMZ1aYnetHOLr+ZcBXTsgWJbLq4uTfLIlcN7JnH+O9SImVaWyjlCPEpIpmp3zpW48rVj
zfohr8UosSWnpJ0cR/7GaANl9mme+c+xXZ2WCqUw9AOQIoo5+TrMNIh6C1Vll9ajLscfhDo3pCot
irPnz8gk5mYRj57BJji5aK45WOg8G4/d7BNJkxIdz2gyxG/mPfjL+jgup9lW+b16cnATDwnaBcv4
EdihT8+L3mOMzw8GB9QSu8TS1GAoeHOIPTtnBFiGWMeRMFg77Ph0K2LLXWgag42QHdRI4EA7yFGA
0ku/JIcyJMTZHRYwXwZKMwaNWgWIZ8RaoF6VTeA/CWBYQaRX1BQi1LuF1WhqlAO3T2gjineVV6TX
RB1INUcKZjIfkMlh7NaO/0qOXuniNeW62CiVtW9UXomQ0vOHb6yHyo/WeG1Ega437waRC77yPnAk
mOpbg02CtK5X9r6PdXvEYEpvFV8R3tIArhM36X7C7HXbTt7o2XRrE5XOmONqhR7Q4U/N5s5gtIex
7XTLlZeSSPpv5tEbjyoDEOaemnLK69PoirOmG+CKSPFgc5hB1T2Dia/GxxB0LtlEOf7RwCQWYbST
lgRIjTGEtt/01iyA7kxC/UmFtqEDOLstr7G1GxX8TnQI5TA/bgFHGltFMHNa6mqp0n5D5hsCt4ar
5ODItJa69iEZxiVcPIqbrORu/C//fXeIOmfGHJ74KYX3HoxafWEZ6UmmGW2kQF2tK370lTN3Ms4Z
ipwYmp1moyJkjRwepx1CQ7mDKsiYpdLFeI4nA5wmEqQ8ZBX4pFjCI6ELL34uNvaMXUiX4YDZL5Dr
GOS1KgDFXcgEBy/cPIHIrKu1CZl73OJuwV65dsQtcwUyYfckowOUriSfcfnGWRFQdcbPcz0BdSyP
VXh+8QjCsxHprRV5qpieM3cbKIs+1pMgVyG6zajJG2O5ouDqpu0XtSAueOGp9ngRwRWSWpjrAtXT
XU9COb2CCKKPmPHj14VNxL0gyWBS/q/zJLa0oOvMgRI3tM6GDM3RTqonc1/x8I2mOO9joL9nbGH3
c2bNZp6tBs1Zszb8Gdq1YRZpCqiu8Vmz03Ml79UX548/OTR1O/Aix/jeU+vEXRnGUMzsuZNsPn+o
HMpZ1/Bk/oGa6wLDZW7mH5ZTC1YT2acz2a2tRgA4OIzVkgK53o+bHYwcPWNoXmYFxiBECPD6bLaU
0Fua1XpxnHANrMcR2CzYS4uNdoaRjmDfPhv4bxDWgkyQ2nfBjw9olU7O5nYQ1rqrXVDwigmyJriI
XO5Sl1NmeykQS67cMy9CE8p/79YWCsfm9z8rKpk3ZX4FY75idrMAMIYMq5EyPbD8KrIHmvpvyZ00
0RMxZPvZl9EGrYicqDaWvvWLscTkv6Rgkt/EYkMw4R1S0A29AIxtfvjUw3R99xQNuh0D3PQnviV2
Y100JCZqkBonNlBID+v5F14U6h6bySjWB4ccD6N8LvFE+zAnK4oGejba4RNmxLubhIiyXesGnDyD
R+jxnzrEy6Avv/5K16TgP7W6rga78QYAkGLJ9Gt4Nlm0s3DYxuzS3+DxjGoIuoRVbNlWYLY/htN6
9pGZJjGXsPAKpS9U1aFPPuQA5aMg6vVJ31bkq7NtixV7i1GedP3Rax00AK9RGBfWBKscL9va2dn1
zhslw6wIcTvI4AFwLABqGJ7D96Tu1t1xMwtDlcCew5JIj4N6FqNIZKgoCjaEWRcwbLkHRzdBFKht
utwO5LeB8NPlXJTvS8G/O0K05SGVfz25FLrlTql9iOQ80oIJSBL0AKh1OO1Od+uP+dRLbbjyeixT
fmy+QsfIvDubvEED8+BUetDH4JIBAQCD1AmNzZAeTodH69Xl+LtdetI1gY43cAmGAU4aMNMflz8Y
GfikN1DbRjV9EUot3lykko4PGHgdcx9kbvzAafmxP4392oshBry46ylwJH5fFybqCI9jgTY7bSzn
nS5K1L1XIsUbjvhefrTZWudvIg+DtMSr/NAy/4OufDVWqueiQvmcGMiQLp2H+rKkBP1BcUhRxOfd
GrzWn0Z0Kv4zqWold7hfxDVPSe5qlJFSFysIsfxlOSxIAHojwdCqWVJEXbKmV7sFT0wxxApCNrPz
fT3q/hM82GVzn2yIcs7R/p3c0uPKhHAZVjs5VxPS6dW8eYJ/gvb7Hcmz3itfPuFpUn86X4Cclcp6
2vODaGPqbVFeH1wDRyHEDBji77BxbvZZEcvZM6ulvUwY99OILtpk/ENe+Adyg794ER/0sGQI0esx
1sCwGkKHq06+ZISg1HneTXh39bO4eyv0qu/dNchDNOfu4z6ZLKLeYNWbexKOnHAr6y3/bs4F80IT
lBGvnJR8exMymVEKactL9pAIkHY7kAau7SHCBO6bvGS8oJFuWDFiiuLdLaU2nn6LWsgUVlzhs+mi
DtUiuABAwUxZdL1fjKkQGYQMZRqZkk9s3NqpuoCkSHgnrkk9cV40T1XpFvIbgkxiiJZjBQAkT/8n
kcKP8G8QvQUShiUuvtjQTeqIOh9Gj5p0qwjY9Ba7L2S5YCqxvEOTKW0ehmIKZMlwDzceQcu2xT0b
N/TRkTKStGd72DCTU2cJuu8OWhiViCsKiuFA9ytqJqG3Wm7DDkCU95JrYrWKHwUIBAlybE1k0APg
24nuBbqyrMUgBWrKXslXl/O/bMgS7J/FKhnrhSgwu940RMOp8ell98glDOV9DT7amLvO/S6t+g4o
06YLpzH64w6D+r5+oWjTBRFE6RKEks/ZFrzi6Ipk4xbNgoHm/HC+q5uJ9tDOdSq7ph2bExMk++7Y
IkAZCzdFeYOFH4wFts2jKK2wJ1i+xh8OFrxF/1cFGYy8dJBkhaCEydSrIQHJvlo3qtm5nTuhqkpz
kkA+S3SehX3GjdSmpnOE9VWiW38I5izGESKGzoiFLxJsay36X6W05eComY0WQ1GdKWmOc2/eQQRa
B0kHvOS5xoLD6udOieqIJp1wZ+axPpr1O1exFdYdJvWbvIU+/saY9U//RXbxJyQYBsAW6gyDHhla
O/OdX5X0+1y6cqZfmnBamJg1zT0eMl0oMXpjn0Q1k/hatimiMQfI8seQgjYC4f/psu1qR7G9/Lec
+oo8CB6Z4KCkJAphaOLLctnt4Aem5ZvU1CNo6ia7bexY4raXHCL8jyqgHzqFp1/7faO3yAemimF7
D9DDlrfUYkDG7lo8qinAmKOZXYb+nI+b9hi30z0hLfTuzBQ1gYYf6UPxUFK7yZLf3SvnSmqv0/+z
xqKrIbS5GkFcdvg7KuKU4BBEiw7IX7BD6+9P7zEQsQBcuJkx0cj/pyjW223cVlWDRGZHzq4PBal9
Mm5x2Rafl2QtaExl0L8IqwoS2uwqNXih/T+/ofcNhRiwBzUJr9nkAG3nyiJv8p8mz7hCxOpDpPbS
dre5JFSWbCpqXWXpEAKTb7iFBItDWTWuioeZKnsuE52tP+mYz2VtqZUYJ/D8fga1QRz45YOMiozp
xvAjaVuyKzr+mEcOnwo/QPkGd7b3VqUD6rSu58FvCq2Zx9k3KSRS+kvf7kRF6hW1kit4VRoruO6o
Re6Y+gIsiCWJS8IJoacI7kC91zdqT9c2tYkugQz4lZI7VPWyd8q24BxZ50NrPQSC/QSKkg0Dd1hm
AVgrMauamzINjiHpdRuHov+l5qZG2XEnpR92kJ6RsLNMqLvV2VOKUh070FYPkThw61gjUWHv4PCG
PftM4GpwkSRWvPg8VSAJMRFv6PY1z5BiAq3OKxYKaMWQWeKFVPBjolQN140oVJTeuMf56aIZ6Yqw
9qfXtRoDpwfXxUm734Bsi3XKoHWvYAYqx6T2Po3bbabFRPo1EowXw5keocpB/a1swmcOSPdX993T
wR16XJUxYm67MYYwoN8vI3C+NUFY95g+2DF/MvGKBNUd6JP/2Y4yZoO9aiu9U64beXfcEmxH25oI
Eb13F583ib39D9WntNfbRxCNZz/3zYEnG/kh9WZDylmrsCHp+J0eXJvMV3PYydGZkPXYCnIr7+nt
ng2PtdJ0ifIpGASspeg9VgzBDLy2XhLKp8Ceyy+IGcF3lhytU5Nh/y/WE53aWmSL0KUXBfAZ6vrC
xxVdgMVJQhBBmQRohGWyXEnpwG9m8hTk+dwg2iGP2acjkjmKoEb9zimqhMDIIQOooh0mT3KDzAcg
BWSvzC5BN1JemEUg5l0To0Y5xn7PdZBHeOg5T3XwujYFFsdlcEV2u5OZW0/IkstSQyUY0E5USR1T
AaZuD6Jm7aWestrn/tG+yTf48eamW237uFQPqw2AvXXOFBQFT9lixTbt/WH3tXv2CfBIX5ekpNw5
GkMLqvgX4Q2aUZn726l+nPuEZvIdCcb21nj0COuKkhKgRSzGU1/8M22ZGM5165v6EiYiiFV9lrT+
gZ8NeNIDUhkMsR6aF5J9Re/mycEqSuBbpQ8uplp7evWXKliO13OoCeRArbetmg+sXUxUg2+FB2ii
qe2glsJKGkiNiO0UR01KYrR9yTk5n2vpjSg5fS5IGchbOSEztCU025KYNzdv7VlnHIRnNf+ctN1P
jhMy1c/H+MRjDNvceyoUmgO6SEgW0ttp3d7Q4C5dBqAAyESawPN+0jLTPRi8KUFmNXg5Gp7cAdac
3lv3IsqExWrZfxMu0kzCU0CKT71nThajHjhI/yZr9XX0A6SCSO9R4OpYpO1m1PugN1/uVo9Vyffk
1Vh5paH+so+4mxaoe2RKt4dwpsvdeiGge2MREpSivqd+rGFFyZ+tL86zFjIRlA1/7LnPPCwIEN+0
99hRygqmCRo9WqA3DmQYgAfHyEvFJJ3O+IQhho8Ccblw9rn0zkUW/13xI3qDyK1WRkQV025JqsA+
xNFaLVE6z4aAiK5zJovHfs11uFWfvAw1FZNQIkaMgL1RYwn5ffsyxv7Owgxpt/tdnSyu/3eEogx/
uEGJ8j8FXAAn1fBnWQUEOX+xUsDsYQvJK5vo4UQ1pcLLYqU9pcLH7z0o7TvcsyFwIPrpsl3HxvN/
kNe3qY73TirzaoT46ASsAYAnrdmRnkdh/K5D+qDvSLa5kKv8jiH/OogHl3F1z0CMP5AtnWsM2yFd
b2BgwUNyETjrBsQROj6x8idEare/NMYGTFE2oCvTkC2V6QGqOqDxzH89n+1u1xFmRYN1r20A0ALf
2/kWPvtnCC8NfHw6EHJ8sALdrsicDNfp2Q7hIN3l9X6F2JhEq/R0uF6zLuHtL9TqJVJshuOFdDbm
ooCIdisIYziiEIWnXaU0xlYVc9Nac7Bi92lM119tPAZ8r+47QrQ4rn0RGQsr/JWfYVfxlBkOaRps
a4Fjl/8Ri+UUwzu9F1aHO+hq4Z0k2Jpo2z1THad4bMhCEsoVq3dZEdIUM08J6mgGre2G2OGyovC0
ftdlJPOPsIQbJc2V2sdFAa+pNKsggpo/B0gmHDL4cLHl5Zb2xlyMBeEZbhAKUVR1IDARZSi15f8E
4Sq8OnoW7AJdi6L5x7LQDNUyoELWFXuqlYKe7xzyUfZgfLCMHUdKXOXnKN2+TUDiItlq4Z4ZMfoA
0ZgSjYmm/u9CsTbxSTpByohm2eVZejay/PSrjenLKSddBlVX9tA8GZBByVHAvxYNfzOhP3yC6e8p
APO+pXfv2vUCg60mHwej5Hq4UPp+ovGtmTdTdCVmAeJF/fYweq+VI0XQ0bDpvHX2Ub6/4Mk5POyU
Qyhc1Cx0+PIP/5DnD/tKhw1vQqwaTaamEGHTu22Wz7NC8XhP46CMTabYXqMUME+ueDGS9K6Y8oyo
TE0o8I22VQxtHKT0bRFo3452+tlw6z4g60WY4CPQF+h4q+CE7WU+dAyGPtbmwqlIciG5hctz5OQq
SSO4I5NOBpMv3qkxYsAMVM7lZSMOG9HPZ655DewxBV0i5JJPuOWezqHUXBNtuhtfFLxuZUkg4RA2
wKBuKU2cJvzXo1O8fo8nAdOvdUpTesldm9UBv7MuZLCEBJHAkMWI1Dv0PTDfvqF5BPIIgb9O+Qxl
cqQQM2+a5yHjrarjIzI9A/ZDYNeB+xAOEhHGwQpKR/0jAf2eofwzUqVE07GwPZ14KBtlhYG6Tcy9
Wa/s45DEcu0XHMNsN0JWDUJKBJufTNRK+q3gcJSM3ye1aFWZnQYJq/ZEJdi7LyyAnXe2TpFEmm8L
DvsydN1qRE63ebKh51RgSkarM645/yKWLH91k7mx6SQjg5ipOxvKSD+Rffn90I9OjuETgnS+Peh8
Nhe7iYVdqWfXNd/ntD7OuUakazRjrSjCZ/ZGV1wQuumAOtKI01gbmHyCoQaDxRNozifVZZnT8gmv
d5BlFdsyWQE1QVX1PRp8DeRxUa7PfGxEz0hGwoqEORo+kjbbLsgI/7stycESzG+XUiXG9DFBakWR
JqZOA4ExI2xLbaYvmY59rHhb4US5ND7KnJPmqZPqhcFhdlELAzLqgKI/CZnrWLvq/f7Ano2bsH42
u9tBqqvArZP2apWxOWOANeG4TceJ74s9sIU1Rm/d/YPRsXEo9cDXkoUg0zi4T5ulxgv5wsKqqpef
xOD4bZ+q5fQDDNYzaozuaubkg6KvOu/Pc8bw8AsNGBwU1kgKFsNE+ibDYUBWbggV6QQ7C2hP5hWb
Gv0bz7bqOOtdhX55hWIdrA4F2vgmZ5hElUKT4IEY5yw78nM2SZrmbIMaXMgRVuZXCs8XjYnWxiZo
reCwG8L4uA/Cp4YhOL81s8hrSdePbfceqvW1d3f8ygr8fsJ3IISyV4gmqKLBjRk/Aj2Q4LW4EtqU
90HK2hniXgwR7VTiNTFon+UqAIdzWlYiU5yDs3JFc5UmJkrHsufO4FEJWh8TnkkexWCARYflMXRb
8+nSfWPIhxn5xwj14NWyz8DZ7n7fOL/NHNkgXZ8+D76W/FApluDMae8UtToXI03w69MmPDoeP0y3
56gOC7CHWj5BTMmLdJjmdSxPGwjsYMO4tG0LsP6IVKZ4jxQIvYxpj5IWnosQ3/ZyKI2uuQEIti/6
I0TstraywF/QoGsfgHiYqxTHiuJ9UwftmP3Elh6BEKtzaLubA1pJPRZtU2A9dtJ3Ruvec01uwRpe
49YJZZyxtvvJpq4je9tJsPyLgVAoHHKOE+KLJB0r+MJCN9uQPCk0wySgMc/H/moYf8FneY6cyKFy
QVvwM83pIIWJf7yDdG5Wu0AoQNy5HrfZeeKrNhryk0yIKcBNISleMTZQTnMxRgbfDJf0YD6T/hzG
BvQYJffw7UMsUcjXl1ziHp+YK36iLkN9CQJ+MtrewGpnShKbdyYsUf3qaeKmq6yChvdbCw4qKIsn
Fe/OEKmlARsJkpya9uce2sv7svBAZrBYR4dJywqtdO46mWa2VyKd2/i4RbRniuWylu73v2bHlafP
8CTt3LtADSktl1ctd3V1MI7xnP8llC9C7W7YUKTVAzGXB4hxrJiDkQz0JFIrvjSdhvMlprN/mrl5
93yf2g6yk9dOoV+T0OgTsJutIiSXfYW61UMc1mGwq16MI2BD+lMrP6J81l0CIQ2xvJM2IUcDDaVk
++zOWaBVA6nAC8rQiLVGor/gxEcMtCOqNIXE97TOtbt/tyUrAKrRS/cZB85wmWow249MBR/aPVwh
ZsBhrqZuiMSrTwC7pVLoHsU8X0zbIsG4WXbNXbqsDdbpuWLemX9pdXRI3aN0WeFWiJ7OihzYCgga
6TcO9TYdDKX3E4/ct3GnvDpy7yl7hHG9369scujJEXCKwXW2yQZs1BUYagd3wY0iy5bkmQo5XqLs
+G6nqhBsg3wFbolIsM7X1dD0t/da1es0VIEVI4QnZHlZDmxY34kFhi0o2TIbLooZiBeq8xKL8fhJ
RqdqI5QF5Du+K8DTTYi8fXrAfGEVnkO6L5XpuXhXhqa+PflsvOmbq8AsChMa5FdCrbwOv5gzXu0E
0tdXVAYJAtirLH5ZFvW4FHzZBt6M3GRRNwgqu6aD+uJ5LBHSvBySHUg7H5lXN0B6IDxSwocJx1zX
QfNajvqITB7A9G54d5XJY8TdZiCn3u5QsgMpJftwGEn0N+TFesbj5+8l3Gf9MQ5mGoRFZKa7EuIU
CmDSO9POnPXEEviAtdPfJBacClO7qTKZ+0sZm4MqDA2/k1UKve2zmS0rqs41s7LK2MLZiiQkj6ar
cW81QpmyyaJj3hnUUD+F6ea1Vt0zniVTxGOeeaCD2cqzV1RH+KTT2IGmy7V7yYmve6w+nQZcv9Iv
Ct6gnMnydt62UQLu2Wav/SGsTlr5jLCBfC2100dOT2B/FgvJrCBDN97dUOH6OMPlfg4Qb7HCnPM2
HVBji7E/RUEh30WtG8RtNZ8cfWZMF+oOuXSM+7nycf2bpHVzL3HVXx57oOEX5F2SptBftBzqgrg9
HgFeq0lYOE6aD/t0C4sCRTVYyZfdjZKQ+536u9zMxUidbyUROn0g7nRIoH3VQL39cutFEu31TdZ7
2MDXWDYy7LR5EoLKucF7LJC8q8wGThwCTYqHyn7A1xTomWcUy2JLlCcAntVsC+PquWirrRZyOfo0
1k/BcsA6aYI5edkDVDu77lrXfJw6egA5qk6yau+W+e/S6jbF7qXMW0IZdo8nDNfvBRReCOUUV++a
zthighWj+TDW7exeBR0XJ143HduaPkCMu3IbhlKbbq87L8X67g3vJer1GChLuQUL71hlxylCIGX4
a/vPCS18V4DBUHlSeu/9Am0K/yvuZ0XIJksR0ahDEBVlOmUFPZE5faP3t99fPpMHwszcJglktytJ
TsJ5hFxW3Hyiv5MzWa3TFkH73FgiM+20C+xKNBCNKJqybu8hN/zE8Dt6ySwWb8y9b9mr/hQEXRcy
kXJtIwyV7MlLPxIXxUa7gBBILw702cm0afRyYqS2l049BTjaVXqBZxeua9+GtBgvm5SGcp/s2luU
ON/GMkUmYMXqKhLLzRNbEr1ECqp4HVOVpeYiVIGTFLYX3wJTsyDnPklgaAiKbHh6PpJtKx5s3pzJ
jdmq2BD45DZ7xf5ZeqbcMe82Fvb5V7vzSfflEi20P2ic1gqsWOfq1htcfBJQqBzfMRjcWGdyDVBa
njW9slSoJ9UqeSL6523/707/Ajzun2lQAqNjRffYtOi87/blmAn4KDO4rVohkUKRHTwhv500eFNX
h9ocFw38FPn8Pr6Y15iWzqMBcndHQpWdjZsyX2uvRApG3jxUrP7wSD0G1h1vsSX8Y5MGy+T4FWYU
KUCUOHaw2/DbbHOcECGIldkAi+boI8nyhgeC3vg388arF61QZa2gQXYzoyMBhtGD5/6egp9jjs8O
gjGmobszOq67Szcj0vYC1KTjvOkmpcR8a7nc5iBVTVrBms8Y/0oa4HOMhZlBOAJt5sIz7igiSO82
uiM5GYUlcZ6Tyk5t0AUIKXiDG7fOlsGS19SjnoewowCyk7jxsNZ3BtW08mBL8h0ARv0CB/ZDfQP0
uKL8WItN6bxhhS1IUXq3zju5VPXV1A5nVFai/ZkzAejww+mz8g/QH8bX2ZLoV/DzmJJFHLO56M1a
N4Zn3Q5Yr4R6Cbe4tw0TUhgJ+dmY/Vw1/+xR6G/M+VCj8ynPfCSVJE3TdFqTT+opE9iWBa10BhbX
mHzYWY3x0wcaGFKuNTLsM4cEzkJsglzs7u3WjdePU7I3x0VsIegSNtqZQXkn6eLZH1s0ok0BKP1C
WfY4Gq+WL2lLICthHWlOO6x8ZyQtw/D8ZWOyqLwcnvujFEG8gegbMggZS7rvy4V83vjawyQFsmAf
bUlLRqMqiOkyPh7hioc90mWfXaGo8FV7DAcNcjoIBEL1wOceib/CBAsamWXs/CTIzkC/M/oCaG7X
DarI13OC4CA4P6G8yfOwawMpMspKUxWhnl1PhfmtN0YOv/LBjlO8AT7o4CazkBHvs0cRIV0jlwn0
uRVDmDKzCu+TGoPzoRDIkFIjAqul90n8/ajQLB98130S67kGDvYkew933g6ag0nc6xh1cI0nYkRg
5foZ6Ap928qoHPiYCGMN3om4VbWBRwMXJkiTT7zT1NLmXSlXbP8Y1WXNQrSqFKbk5fpOVgbiTanJ
H1EGTSlLoPeIgD5/iS349xYBplgGSHB/ebi9/zK+jc23yRQMiZ3uweGNHk1ga4wTGZQwOsBE6+tB
SBCDE72IFiBAWCrbcVs1Bs5sUrAuIDhGbDjgirNM0LW/FyMzdpUaq1aBZlVm1/F10RiiZApYhmOa
HwbVO9egPUrz/jKQ9tbSPnAh7WDJV9sxvBKiQkoxDMfo+gCrYyAeC9VeEKI9HcQ6H87PyUxtd5IE
4HDI7XUT9kogJRbM5D2i2TpuKb1VYQsQvRgRxkpgTTKf4nPA7KuHFYuD+UK80Wx0e0GyPQ0amlGq
XIzFotvgF2IPBG4n4QA5H86ZNg5Z8EgLbop8ZxU8gWpQuRdm2BObam5clv+ZTnbGViT30IYGsieN
T6AOzM8VtkPXBjen2WdBtoCWRH/2wYfK5L6zkb2+wNoASaR2ABmXVFOJ3ZdXm46c4GHfHmYXPbNa
vdoRsxLhhhlZ3E6pHGZjM7R/POXTbaJaISrzsFQHkZm5wxbzoA2XGQGLeNS13TLWIsm6VKoY57GS
TbP6S4GFrF2CVudWVHKCfWMHBOAjyN6w4+tjzQYl41Pf61N70UBEr75Gls2gS+2K1I9NFZkun/mx
acgEcAWru4KMXqWyoGz1hOnMwMv0nQaklMO0QbSkLSxr/x836qExdxeXlBECj9DZMx5QaWmeiiNK
a0tVNTdIF4Sn75qIDupYvnf5q0qRTF5jPKHzjVsiPOLQOnJQHNtgvzhMhxopV/Lsg/uRHqbVP2v4
7JRf0MRDm5tiGOjSpfkH52Qrv6Ek+I93iZ+XSelJ9l2In0QnBlD31nvSgcjpbG0UMTHXeuYoYz9G
ZDcW84rddHQA/Ojyf5SR9HCYxVEPXDDjmvazBSKowsx+2SKesTm2Udz3qQ2lBwJ1hbZguy1M+Fm/
vF1Lm1yRNp6LjVyX8rjK1FHxXqy6Rmn+1hV/pYl95GSM/wOMyLL8pa2vKCF3Wbt13OVQpLyMOBCC
WhztgQBO+VmBjkpaoaNIiTOLIZrOlq7WuBeoCn6xSdxQz0Wo7CqFsYeJiwlN0bV1z6UZLzWLFtZt
GzmJqvFSoOvDM+ekSAgjrkLWUAVpt76LptOHbcZa1cf1lw4f+il7VVV4S2p7qotUiJo+28k+8QPh
1toumLCAVZqTaercY6bB1B5cZRkzlCzaE8B/MbzMFDyrlfAnncEp/OapwbJv3oQhgvouh270kp3h
t3e20uR0SO2b4Rej48lV5WQOuyIQhoGvGxj8oHKRiM4muKtsOzM0O+OAgjK566FL37ugPZ3HvA/5
l05Oqc+nFIE9bg304oP/w3yANkdh3MzIUEy3YiXM6flinedjw5QgoDSsSfldqFrGrdq9g5CQ1aPn
tse989VEJadq67QTZkFwPLDewyg78f3l3C8lDn/BJ//J7YzP37umXdLLPyVPpbcQQHXi/qYltGXN
iEWIeNDjLOSLIxEjdo0hHvfv3BKxvQbQ4HCFlyRogQu18q9EDdnWWAEHWaXCgh+cjk7JRp2Jhqb1
bQVuHh8bNo9//ohYtwNo/sxjK6V8TCdkclTUTBAnnvM+od50oRJNT8Icj+NkJm+8D1f6bbmr+2r+
L3ode8Y9pKWE3M4OVpzHWgbpYPNl8xmLXbUT0KH7dOAKMoKvyhKFNmBOIr5LqRvLqioAAXNafFOc
rOixM/Gaal4Hz65NQ60PRT9pvNActbAhJ/oy8xz5jVhQlUxqYr5xquhxbR3CVDqIhhHLn1iyormE
Dmdoh98pk4IjRAElqtDzoBSK9j+/fiQsjdf/1XR72mm0vhor2STVAbFwxxusVWdmQMtmqG40Pwgs
pUmVuKK7iNSMlk7SUhMnRwFD9TiDXiddeiNqXLkpVAAuJfMcgvn1lgh5VPNrNLV2x6EW6QEl5FUB
fi5bZ2qwQ4ZLXtrLK6oSuZH37lY+NJu9GLjBZvhQBZ6asg46/MtKds2He+K0SdGgq2KWhOB/VuVn
TW//qQM0VIEXHTzPo2Bk5CpmLqTOh1i9qQiiKx/blb8PcP1sOUoAO7fBz/4hozeMWqtzF2LVV6lS
jVyOGWqMBaep4E/K2kRrpwEoaFUJkMzE7GCpIcy9C+DjoGL0ec82mT18ZzyfiQLUc+U+hMMxbIUT
DHd2sUqJpHAzHEUyOHfj2KF34/73qcqF0wr8HDFRZEuV16buqInUeC/VZE/eU18o3Ga2iLg4kid5
hsGVNUaoDlh2aPnelmEYAe/uJpOhhhBCDng1APhnyJgsDJvhwutn4jppuA6K29cpPKm6DQKTmyLr
HMQWLzc6nqC/Tp/AaoK2Kn76XmL9s1/Rf7wUIytVeg/6LeRAQWsDDxMne7j1eFHMgc6N/ZmHl+H8
4b5ewxZakjB7DeooTPrF6S+TbzlbokXZW1W6moIBCSA/kA51yHI5HMqJvdjniiGYNA/ZfWMw0fir
KOidk6/9e2nTkQS3ts0u/XOxQq21CE27m0EZkKz4suSBqF98FMOHt4b6zCqCno7mkfMb4JVe5bQI
LUyalz/sgZi+jPFfaqJ9nXtC+eVGIL7nnq5f8RXu00YN65bdfB0F4agXt9vQxGW8gBBbboeL7eNs
cLoa6KlpNT5+6/TzsUeE1nuf2qNYsDvSPBngF+Mks5nVdhnbHZta7utdspL4h5yH6T+IdBcZYPNY
nPo5wooXjIlcPtMVkhGeEunHC+7SWaZOvL3bn5+Lo8WrS782LYGKE7+3reJEuDGWFR/areNRuE3t
hD4ZcV4rIEi1RfGqbSmkGIyBiTJJl4ITpE1pdYDCX4wqzliB0icdT/qgivjYWt7F2N7Tp6kg0xJ5
18pULrNsofhck3wxkyuwpyfajJGjmNDkNjJb1B+9U6HygLwp6WZZIoM7adwA9NEc9ZHx5H8f1qfL
DGQfGMyiF0eax8QTxm5B+RoVUV4r36haBqKhYPaNwGc0zAOGMrXprOtfIQ5DqqSYGtVcYTLn71j2
D3BNrwScR8/2+pnCB+mhhVtlkO0axILixPpS32TcYMmSd/+T5wmePz0lP8RwXyaSLKDPCfr8kZYv
LqvMPRP6DdxGVoUcQbXGsKO8s6AYuOMoo2pCL9wvHi1WhBm3gkzN6URab+kqBOQzQEBA3XVcQJFl
tL1sLaf94dskczr+rrY/Co6TqULLYVVdOuA7JaoIRpLcltbmoLihxtVRhVXPErUA3j9OsSmxDnB+
ddgkgkBe0BmvGqUTrqX8Bh5US/boE5ku8OAnf1ujPuV94iKKdPlA6NEP43jIxapC3U0HzLUwg/Zr
O8k6VP+13pSOHlQ14Jl44D1ttjQeFkfnBAxy1ns8oCSsvWtY/z4nXBj5bvuE1Xn2sG7lBLx6WzhV
QxWZItoMzPkaP2CLi19Og0Dc3mfPkqkYAbPUYH6S6LR1nHiJYL78Iq4e6wM9EGdQky1uVXZWqfwr
HUCCOot/dX3dJtZrXIbebHdfk2vOqrzgshc5qFpkcYVAKrEWPFEX6tt+nDfwWD2phzd9LgNSQZtF
AU4AMxweki56bWFDG23yFRwCZaRq1MuUNy0WEEyDbZzAGJfQvByiVUPQGLA41NYi5NfoVwtQEXdS
7uaob/DXFPEDGyNCvDg6WXgYtvtqudfMfEM4KIgc4dRVSG7d5U7h0nrGEmFedVDjESh0F5XV2Tbi
RCSx1ly5lQDMcEl4HJgeZLO/3IZYQxEOfTPoWIB0uCL2eKHS12rVE7zFKN5O+WM0Hk5iFS+EdE6i
WWLagQ3WQYY0QF6Em9B9a+q+VSsQyIxcHR9CqiigexXUGB/sB1XX3W6GXsz9flh3JzLozIbWy0fp
/9nTlz0w4U0cNiR9DVtlXXOwZknlFAIFC86RhzNoxWv7n4kz10toCsKYv2RRnaHVzvQevebYH+ZA
Ix05Kys6rsudccmLrGutncjuejwaZOFuCgJMMnNLbsgb1FtdtEnSuxJmABs1JUJuMBFlNXUQJW0V
HU2OIVitQpewdcd7qlDfQ+9DR9gJNSPohioheb+BC3PBjqIzTMgbevic5O1ojOsk/1cxTHVIQi64
/00syJ515CDLKOYS/CZ7z7OFJMwVb8esc96BbrSlRGz5eb1gmx738IZUf/M2CEN17zY3pCRGPP2W
DVPYDag65QbZC2scDDlGROEUKIfDY+BatucUvULDY1QdsUBLkscN3HmKB0+qrsk7yJcpOXmsREN+
DP2awxt3Fvl0JFv5+KadU/Tp6es13chUfa4/ukqI4UbP3NzEwccdB+nv905Ci3bk0tU9aC2ETDFu
0qkZYuRY4e2cC8mCxlWu7i5YqH/vl11qON7mCSNgUefzyPVBpjB0v/wd8+v0q1ahROKSUnoHJ9Cp
KMF+TqIPMcHrwbAD3BdCYw7ozrkEdL0Nby6njwYbnhzDSlYirvNMYVa3AKOSbSfem7Y4Lo/t80Z7
aZcpXocFhw2N+4vuzAPJJmmeHEp7IEqmXm1qpCyuoBACIjLcfoPq0BgbbXdPDxKNekG7cVR3vcgi
8LYiCdq4LHDaDfGCWRR3BDafX+xEzy/UaVhwG+1t5oov7B8QnyHXYwt4a58+wmXoiRAEghF/GFro
slANYoS8Nqkla5ZiIbI/LOJ6n1IFXjnLFpKBRJFf2d+E9/vZDoQztqt7JMZTVLudO8jFbm9IoYLG
kAU6QVyL/2URQELKZhEHqfsCtQvQpCZ1IVS43oLHf0I9wTlsOqbdJxFEMq60iqoc8FVnjVkd1y7X
IiLeON7/hHN9OQ9j7kuUdpjxQ6Q+7cazihnzE8Z3r6vZwEx8JVMxJf4bCR0QjsYf3oHuS+aMQhDE
SHptd7YfPbAHSLs28pF9pCu9cqAcE6RRmpmLD1wfn2Hij5KCep361WfgC0bTq1o+PN11In+bpCjj
qlavaPYtcU3FAkLeI8hy67Tj3+iHGWTqXUFL6G0ZVnATgbGwQ1SrFvAEVz59+1ltfrteqSaLZz+T
0AB9aNeviYKQ5AtOmW6uIzKHYEuKlEBVYnFHcoxZN+/zvuZL/XR8EbXhfWjL2w32uwxV2f5/BO9A
oZsj7vMawvOJLac7HSKNJ/hqCE1aorUCChY3pX507uLP10MZz+kNsz+woQ9xsh8YqQFUzFWVuHrE
lFtoLzpYbwlkBpuT+V0li6xDWZf9nTrEFajTiVRPTdRJvj/RfeDUt0TPlbLdB8mhPluz8th9VrNS
1cB1I45480egop5m16Op7iKQ7BScKrZaz1STL1ipMBqJ3M7XZbbqeaqZaDNzpYzqdVkNXGI0rpe3
1WPZ/7/hFY3Q1/d5ee4hkjBTXsqK0nl+xK4fKziMKJ0EsPN6R2EFNgbfGmZHDaBgIYgJLr+6+bZ3
GgU3ZpUIEY3USPK12NfZJE6w7Fqg3H2EW3lGTkbcUwviT+JoB0qaOR45l3GiRB9ttDKaUrAmTtBG
yv28R6Eehv6DOtN8Gvyj+MMZB6AiFKSaF9RPJHOVn0TN55n+5Hq/uwzjajSbStpZdcYj7MkuNMSx
BgsmgAjXi6V2zG1H8/+vnpY64CAje7z4Z0xm6+BdYWTz7RZaMCQP+6nYBFHji8uSMRPwzhBfs93i
ZBBCcZHitYw6LLV11m1YWuEWp3S93ffkH0Tln+X8Ayd5S4YHQ842vaTXAswk+Jy2tIz+dOiJMsUQ
xak2WRqcB4GJ09p2okX5ZzwB8rGZws0lDhvi8KiRoTDWTIKKfwZHwI+oyD1W9BqJqK5YK8zETeq2
OYMcH5SucUQ8KAS7Vwd5D0WOkiELBC4kHh2UTQ0Mgh3QyrqbSkXv6nZjv/YKpDm4V+e4Hn9TxELk
JKSWgtRPcZGGKzihQtQQ5CqUyrIn/lXxA2W7i0evvCmQs9JsrjscwfJq2Pw6leGWIKZPlsn5hD5f
Jaj51cqKEd+DkUCrwILGbdKSqEl6LM4qmPP/jWGhNgfULMPSWPN17wHVEjYDt6wJe+1oOr3/7mZT
vNqKWgdeCRf3da4Wq7lPeG8n3TpQ6RwEH6/W6xYWrUxm865Jj17APQrwnrQg04C09wl7Q+EUsfIH
Weu9+JFKzfvFT6qmvQccI18Si/ooooJZTL1dLR6FJWsRZCLzN0kF3/qdq+f+7cp5QvQAZlJpn6V0
qhecFCiVZif5OSRWR3tFJ6mOX9eqv4aDeEZR4kfZU2wpLUF2L9/9puLBJXove67NhZZRiLOvM8S4
Y9UqBiXJXsUOSxQdgBcXZYcZksfl+LgQlOooIRZRDD6MY6TGfvHinn48x46ZEDQAV+gpxxcabp0/
IiL0wGR+ihhgnPZ6+A2C1Q91TNr/5VlLn0AqH/tfQ9Q+fjm7+KVQiGCm46lzEnzhf55oh2ZSoRim
5M5gsx2/tW4Mo07l8w+NDWLYXr4S24nfEErTXc3mCpZ2Ur2wadzu7OxzLatV5Fb5ZJf9o4pgnAL2
yWAIjFnnXBWYbaM7sPXj8KdKEHOQ01teqDS5XExPISgbZuma979Xa2tUBq/c51EdPeliohPYDEJQ
zicMvoG/dBxMv2sZ+IEC9JergLKTj/SzY7UCLnik1ZNI6Gr6AyuOjE1tVPFsR9Q/gNFRtEzTnuWQ
RqqFTp7ZnJsNsw2MLrkiyNe0cXKYomMeaqpNC0HCRa1mdOaqXWY+wPPTU+pD6xV2foJ1C1Fay8JQ
fkofANccZVG72SHZ8pcIiAp5LYDPYxvLXnkZ0IV/0snatzqUKXvM2Ozd5803MMJB/opBwZVrZzaj
AhHAusu+UE7zfjW7/55Wa+PkCV/Tvp309lSsBDsJRZ4lY1aZAu/mbcirC6aiy35AGJ/or4JcI1vo
d99dggmHvMzXMNNaaoNvfOKGkI/VG92WkTzy6s4zHAVzjK9aYfylKJm+7egIHO+VYcBKbqqnSj7e
cbqXVxy9q6YbVPjZ9qZoH8F4bJfua4Zo44crUUptB4YinX4EEm7YKFXIMbnsM9CGACUmExz7Rl4T
YHsEUZUFwSvK0LCRDYziorSnfsfQl2wyY7wn70e5RQWPzwcyytX5IBNzoCq4C+7cq8oKPEf4SHWf
MwDSMtVHneP3EJx6ucjLetQg3Ww+m+iWPfyY01ZNIN3XYQ0anKH6KE478iPuNjD2ZuVs+c0hLuhM
lYXcx+j5xj1BNu5/1X8lPWokThGDaV5w7JffBBXW41BMJ3n6r7oJFb8krFgA0IrV261q801ADpaG
yFqVa0mvjtSdUI/yt/NXA7lxMEZcskl2mWQwqB4IP+BpX/aS+OAlzxdCzuhK0Hq7SM0i/svxDlVs
Ktmt+exo62q0zX8bAttGcqFnHW+DOR772vwPymSt6PP4CQY+buawK9EtnjihB4AdZGtBhabrfD+c
78bjAH/Id4Qa4peEVcEIpzdVBW6YQUdZD6JpYS3jbvp63P044RqkWYp22Dsbpp6z9fbwyCnxL8ch
4Z/8aA8mheOrLpl6zpYp4EwDCIu46kyd+/0TOlsAc6kn8Xg4ruVq/arA934mrbJf+HMipZe+JQV3
/Nd/e6H8EFGMer1uaEL17s6Mk/+DsiqiAR8DdhtQSCNqpovIkvkffXTDXAnVsk4uCWq1oFZOfcGs
i5Qpq0mmuDP/pTEHAW3EntAZCsWqy8kAqKTiuBgdoMsHDKy/D9O7Fm7oiASYsengBmZtVDS8cG+N
NJ6HZVT8c5KnSJEm/Q3fhrL89oxDqKNZZnUGvKKH0Y4jhg4FPzST3bij6yzfA+ggAvCN/X/P+cag
hygBO2yxmMvROIDpwrNdjdNpVxVOvk00VmzjfTTgNMYbCGUOP+59IYiv2lNzFJbA7Yj3/01n4tdY
yqRtjqvf2/0dDl5pNQqbdoL2YfU5e/qq3v3yXv/6xHbwuThJekuv2vlxx0AXPopQCq+yWoo/KMkA
+/u/TsnDRvdD/2/ptnyGwYI16VYiVEZIN2GkKMkwtmX1tI3W6SOYtCbNeN4yiFkV+zB+i8X4Gpt9
pxQ8Lcj6frLI0c+zEkyjmpuTOVudhlI3NngLT9Svga+AxSP6iT6EGRjYytHkjsoORt4UEmvfFUZs
9lMpR+NFfgI4ivUQmctNSrHQTUV/TjcStbnYS9FvsOvL28ndC0X6JvNYeQN67kkhkZmbGnTmMlCs
n8/jenKKZq5f3FJAWpgalj+Y1BkFxXpLWoI3odfxl2BtPtYPQNkJEd1C4SaCgkfzzDol+cEIRDsl
Up6oz/wcvytrK63z9N6tBY3iEea+k7ASafAUrm/PevQx0wGTG5176X1LwMPSJGNUeIL/cTHib46m
IaNv4Ma9tcOwduSxpG7pT5h7BdQ+mXrb4vw2HAeJSWJs4rLYNQf4LPH7fbkYJ0Sui2wAfH72Tzju
GMn9z7n2RR1eYTWFymLXmnjQB6y3AMB9tat208gkFSi1fSRrhbXXNf40hiqgGnE//Roq8/S0ARM6
Nu2W9nsjtvnvR75rW8RltXS6UHnjchCgnVGtf0o+S4IAHJWCuJlVanXnnfBIYVWsiuYajwEYpRx6
6L/ly6gVeRXi6UOUkW7E7J7F5WKXseiq3VfJKvovoasZ2ykcAylT5ZgmXE/6NuHWbvgHXAYdqiOL
yjriui5Dbg2pUEGT1RgD7c+4TDkgeYX3afjgk4+AWsN8aEfg048AAGFP/wG698LFz72bVjAo5kuh
XKt1s0eq3z2EdfCWnsjAGHi+9tgiRdaioiY7TkVGy5TQCTlaAhFRK7jqhwDgOC/1dcJ6hhWg0Gck
QUauIdv8Gn3PywPOngtYfzG0VnI+JaKDvMTfhdxzmgkdtxSgrv45oPa96amQCbzqWWm9sf0KGT9+
tIj1vqhUPZYJVHV0FjROSYJb+pvLuAp+o3amOdAAHRTvG5nxxc6yh2tvMSBGDnaaZ52H4S2q7mgl
SxVdJVse+6jj4RZEj9QqbDatEPV1C9ZN6OkAHWQt7v1qsqB3Zc+FFc/NfbFhmEYBRxfwPfIHmBD/
JwnPbd96HG63GVTlPXNfnDiDHErBYAxY6Tr5UgCnkKvaBIp0BW6wJ6XUuGjk/JCLupmJ9rFvmolG
n2tlCHfl7bRd4RQNlbLnm99Bd4loCIzXD8Dcs5Ku40mDsXAMC1kO6jTArRc3X9ZOrojlDh2i90kT
Qkr5nhqMOWFbXMfJOEjqEqtr8RATBo3L+Cjz4rlluIwUpbfe0Av7V07fFpCit4vbt/swi9LAwdCm
yS7Queirhf3ewGSk/IJuUyfhJi3sWY95S4M2pSPzTMgMcNQxze0U1ml8svhc5n+pDLoe+/PZgQJf
BPOuSNYvIJpFHHsPOviwFenlkE+3UYoRz7EetAAvANT4TjWzmNezImT8++3rWreWT4qpMe+2gBoG
ikKFdorFQ27nJUpAm0Ds2gcURCq86TQibU2h5IBPuENGM4+8El8VJxnS+DgGCTtT/YNU7NhauIyL
FVaki4KVDdrdxPC3Lozp/7lCEIj080pZs/H/vk4K7db6w/V5Iphmti6taxiMEodQrEmv2uq+H2Ak
LN3OJgZfv0GeIDqp2cPl8mHmtC5FfQwZzPNMKxdhNvV1uRZtUFmuqfu3Pc28ebqXLZp9cCsVu4Lj
AQGGVGxy58wVewQCwA19WBQ5fOBuR5eE3VV5XZR3Umlj1feRxpAfzuOiCH69EzjKDX1v3ahZkpsF
xq8n5SBe8owO5FojEurG28MmnHZF0WWkq3lLKzbiuan4RO3HYG6Q7xCRxg6j2iX25aFkbRNTg5gM
5qqKMxRr7xZRd9BrBfKNSNEBfBwKOv8nK4LZ5NIMasCb7+qrRGbl53lGCEJfx9Dj5YKjdT0PgK+O
yg0cgth1sEzBZVEk77AeyhoQdWUfRSI61thZsFLhg5npKmlgtt+HmRTyoPsaLc0UMJ6r0pY/gxdW
/UZtYTEv/u83PQxRz+XcYdw2Dk4BArbdypZa+Fc8eJthDSqY/eWteMNHmFNHT4v+1WLmS2+u9bB9
CCmrnYcTCEY1kqQ0E/YNCBTOQWW6FfNLJ+cNv+o4HEUFV80vfraXuRopAslGSoLPTnwlCk6R2u/T
2SAhNUZITPA3erM4poWIcSMnZTn0R7ojv01uoA1GsNobTHZ8Txb/S8oCipLI+PcZ6tDxSNToeV4e
PN58GbuL5Yg18XJEfSXUhGlNLEdzKxS4h8BPpBwZAwf4CLX+KaJwICYXRRpZjhBOvvYwxvcvCBQw
0lWpdvH+yHomwJpbd79kvXclD9ZjcUy48GyJapNbT39ibv8C22F4gkeml2pQs24ykIm1TKrNQoHT
itAvDet05BIZ9GQTgu/RlSv0pd5UlQT63F3cGE1PWc4qjkZ40c+q2tjPfytTV4Cvrck0bTS3JAAJ
VCYuJ8EHIaLEbTpLW1UahU2WzQ+6f1CyC/0Hieg6HppfORbDzMLRrMdE6FlVwcjPvuIuSnLU3AXr
/4IxGzSNKzmY2KLksveZITGxorBE1Y9ZqZumuPBw+JQhG8UzPzEOzCBrmFafwEteKhrrsyo4eiKj
Wd9eaPfkifk8o9sqbtdoBtqNbf+AHSLmUPwTXxndAosFTuc7MFri4i88sa9ZtzF9RkoRwqILZI/0
zsUG7lzR0GZ9MRKswU4q8HFpbUp7/0Ah1Yyy4yZCgbaUmeBxhnLyTZ/GYdX1ZWGb4c0nHrYFL4NW
co9kgLlWVTmZrn9Plpq8LmwhBr1pSTLyfy5cVaNtsoPVJWPGQqLyjOfecRf3G1V8kzPAryOtwCS/
MwaGw0pWf0ouGhYoNuBm2T1a9SFqecP80gKdINTFH2BMLtcUQvmdJYCunuQ5M282z62ZI6+5UHqb
rwS2i8MiNzcItcy49NJ/Qyb6ePJMipCDpFQOm2g5z4F5WAa6JaaPgCWeStnJYQAFcIzNg0qsiarH
Wv5bJ3HIUzXK+U/wdWM8k5qtLolBNyrug0u2zwfuqMFrBafgUlGdCf8NfnYDqviKJ6Hira2tramU
MLWfzqvIoD9KEJIf6M495upoIHR9DOT3sYmUBNBd+DlqqeVUtPR2G4uVAr1Vch0UYbFBfEvd5NJw
opuRay6mpv1Y6hrkXYPxboHl2oRIWtLoxk3mC4LvQ26iN/xlvDZBpHBh5W+1+E/JHoU9YHWHqy0l
UdMEfDrjowzbR1AVaIuqKt+3lSU+StkOSeHRMlmNDigPZTWPx+hm2MuPZSle8XAZBf9O0CF4uW98
0Cx76xadwu+wt7l051N8EGB99yuwx7VfFGgQegB2WOzcB0wz0UdDVlw9zyr0DzAWppTMk1M8rLK2
/QQmk+2WsU3/uZ7Tb62r8pAQCiw3GbHyCnhR9jAi/rJi8ZU7s7v8lHKDsE/an71x+jRe5rzHx9+n
BVPG5+o7f/hRFOwFunEpqwxYYh09SNpnKYM6sZnCMK/5yILyTf2iBvgqk8v0iSM9TSmqwomnPbWT
fnjSAIvDPiI6sk/DQzwRWlUJn3zctWXDL7HjHYs52LwRzeLag3B14SPK1YbkvGy2s7qYEzIhPPek
3HyZKS1N5guDqqjbaTr08cGPjbvkI15TZIH55L65iCLILwLG79DYQ9Nn2zgRibl3xPCynmgVKcIb
woMWAyha+sxu9EyDfWOtfW5NYVYtY5lDkO32tM2v8xf2KyzZG6WGdpbXDjKtEBHRlOMUjMC9yuij
F5GiEQowy4SyjIs68Rg4YW06SBl3UuqP9Id2hLfnvuPMGGm2pYsywLVAb0ekPgGXPCneyf3i/toM
OadEyl3Cpvwi0xOtZFsKZQWMcfUScou61zgc4Zj2749hh+SPdcwiSXJWp7LSmmwLLBnbqlD99CVZ
rwHN5rMfT7dCj8dS3l1q2EcpVcTLJraRcwGAC3APrbXDV/yvFTrhlpMr8ZAqg0+KrztWP66Y7+TT
/ad2N2joNpM34YdBqfpMhtETs3dmVbcm+cMaRMP3iAY7BZZq55BpAkFSWYKFED6nTtn1JAjT81+c
cRDUgk2PadUc/E7VNkNCO76flfbKK/macqsos2B0cGXg5QhvKUJG89kWK7vEJxG5YWIQyZgJQOQF
hd0muaDvW9+lYa45X9CwAWLNz4W/u+6zP/rU6oEm/CSvgyVhAViNBQXw3K6KwJ1Nl8pDUyuHXVR2
tAeh0sEpUhNgdg5tbfmwZ3yZTMAKkPNXkEvfaPMroJxZV6CzD36Q8VJjw2asp/ndias8JpEKy8PS
VtbD9vKi3bK+th+F36zhfa3/lYDScuKr+xMGd1wUZ03qSxr6zsm0XtFRBrmmKZaQ32zchyVf8ej6
1GtXBoh9x/U2YFbwbBZ30yJgTEuz6dfu4fNQF9EAfMteZZy5wC46z7UyFXXqSFN0aRNcWgxLsV+M
CLbcWwY7QUyEv2crpsB4xCo7Bc4irTuPjdxSZi/PjWWT/Gedr5y3ue5D1llUmPkCLXqPoDR3qMnC
uAp44Jv9jnG7KDn4fyKfhMQiP2NPo51jZSYUoGmZFyNo6nAmgSDGavmp7AgkEvykHB2476cgb+F3
A9VblyccG/F+93txGPLAnx1N96/eqn2oJtEqkQIDpWzlF1n5EZQAEHk0jH8eP/aZgD2BfvfruxHT
1AYk5Iabkr+gl14XsP4SQ9u+M14SFMds3I6tWXFlLDw9zliKYkoYongZayj/QhujbTAzo+vBmgkJ
vbKQs5qVnfDCuDO0YW5QRso/zv1p13VcoosdDti8aJ1+btToYtbboCv76r99zl6oNutrI7NoX+vi
YWU4JxBA/X1X6TxjrmePtj7ZNCuz0hXnzuKp+hzaGnP1erxLp+lovxq60Z9gd1rrd9+3xFqE8P/C
YGXtCRfAIzkmTjPpykRHWZweJZN09IvE0/4cMlTGItv92ue29xVSmbJBhuQEdp48kLD9YjeohQyD
rZPcMwV9264lYVWb8qJyS4W8yGeuoF8HeIw3X0t9OXoVBlJhI2sXUpcBGnt0SeKCIOkL9m5FLl+H
IR4DeVM6d3iKMCVbO/LJa+/y7h8h6jszOklCcD9+sqGsXKLOyhLCOY+SZShbgCu32ixDefeB+1kw
PBs8TWU1Rk5sCOlRcK+mNrsFUdyz1J97xHUxVmT6v24eLVRjo/Qb9/nbsG5v3JAKY7kqDIW8SKjc
wB/wlVkctvByYkru9c8gC8lZzyVFappIM4iJ0bgv4NZ1jOoL0Fa6gp1K4nK20Ji504PcBDwpEtcw
bzEff7l+ULK9AhV0sZXvCLPMa8eoYUfZq06OleFXuntnnTCugYuZmcUtO6nY0yU0hZuvmL6Gb+4I
YQrEEzNJTrRo1orAxp+xhhD7s7Ha61CRLBiTUn8a/jb7wI38oBY+tjDr5ld0jJPbyBWdb/4Hwi+o
D/I/veu4lU8kvqrrd9HqTcHYqqYAvXzOmbuq1jFVIfiAEOy0NgrkZHKJuyedgNhNuDTZKeuGQu35
0X+RQLn2gsBujFvCn7cmIrga6SDK891bkssU2HvY/T7HK6TuWdU1EO5n931PpgzOis0E+rq5N+BG
OS3rfyD4dnYgVeh3AgVH7RHuauAgu8GVcRKmW0S3jdPkqW2SlnSIokZCHjWNWaOM+XTParpIoCZk
6VSC5cCXpPKAEjQDZ9nzj5fOJOVdJIW1pu5Hlz8EhDdahj5emCvlpWzdserOUosjYwzGH0lfmIgt
Ti2Wd9p8V0R1X3cgpCT/w7fDM8WyTM+5Pzlwp/fUnDNT2bZ4e+swF6OIEBUaAwBWq/uy3o/d5Gam
VTv6vvBYN/PvTY61qEpsBTnvr228DLPfYqmSfAWr5UQ9VlswTsLyt0+ZvhR1/3Meh1DwHdlT4NB5
jewYTOPXUXvj4A9taC0gl9HWh/fMEm1NWB7WY2XsBrqgRTYQ/EiOWMRmD6yrL1EQTweegMtFM7rY
oOi2WIJ75IX78L2f6yXbNpl4zTcCc6g1Kw2blp2gTCI+L8TS/Yo0+HqpvDpzimCrpthUPFhYvTQm
XcciGg7YHJx9Gx/yQzb9aqLRdlHYiwme9CpgsNutLoV78kE7RMzlkRJPr2ZjqZ4ryASdP0pfkKrq
v/ewTCDNMcb3a+R6X3rJzQUuCOfcrfPrKlg4bthuyrXdHONY5zgsnUhPgMrlpi+W1rWluMMxkFxw
KnbbeZdM7vhXk2wbYYHOS2vaan9maEgrPgVoatxFnJW93sLnB/HRlScWCcF0FkLEWlWTJVNAd57t
PzS7v/B1e78kU2d38sU8iqhENioSpnLfWUqaXu1rMQymPeNMPdBI3SZ50K57RKmaKnvAsLLtP4/Z
q3UhhD/hEGXhuyljjRGhi/esBCxn0oSZUjgv0MsjEznQe9OgOIS0jdNICOY+n9odml6jgejlFFEJ
Y2XkkWo8HhDzK7TxlAL11CZR0VF3iOyuH8qI45mNArUgYcOSzN9Q2qqxZ/nI/IoitQrzdvTgopX+
cE9vGjIs6mWsCXhZlywjOac2tunNnhcVEBpDHa3RlfJkH6FDaqaU9u2WJauiYYH0uUu+rjfBvizb
VW8P8VwGV97HVNoKGF7lSE9H2GHwEFxfUSlRbFm3Q1MhCKkKiZubb9gkrGrmeBnyUWRDF59ua0hC
aLmzuIqh1zhT60nOPBRDyXvkw/hl26yblNLV6kGf9Bdw7wujWqt3MVMR4RdAe9YFgz9FU6d5NXsj
qdscXa42wBCKwS4yFx/wvXPbXPoKrQ4lYWm6hkUh9MhINMdaGmLsyK10OTqX7Ks8JOaz5AOQrHuY
F1oRNYSFLcOBy0BtcFLsooe9FfYnq+eRMILy6/DL1vPtU5126n45dtsoxNGWnXiGtSxhPtUKc6A4
ZmROXjt7MioWJfMlGNs84K9jMI2SEDJ3E3clCGIUEKYxZ+lfITOWuY4O89ZkUDSisvEYpM4Hy9/2
O8BD37j2TetazMUc1cMMJlsK2WYZDLpeGNdNH17HJXR/zJYrtG2K17P9JKx/tuijgEMorayWvkW2
UDDVdeYZooG5Hm/gq/E/FMCStoXVQNBRfzmFMtjr10kq4WulrBFmTEhzjjGtfxDUP3zwPO4OzTHC
iuw4K/ZWnENAb4GN06H6BtldRnWWdx7FXpaaDrW7z78IMvF+NKib0mFl15UG/SFmKN5SbYAMhovV
jnheGgusxIJNzH1U5bvZd00+1ExUyZaXNNyo45cVV/SbFmpBBzxjimaYyIvHyTANjfMms54IrG0g
pjYeUsp0nAnQZD9fGgRd0s0i56RJ+gKh9V5spn9b/o2RHxt/GVSpp8pDMKD5F6LYF2+hMqCrtP8l
CtnO3mwsc2v3Em4EfFdfaXB1G0oT5UVREdEZlBtOHpnSc3dgIygpiu146f/tFPFXVQuGOXfXjMZO
ArY+zeaIwcSBdYrLiArfNU55gurB81GXzayHPAEnsLrrbHm6BFpHbWy98xbE1jD6oxpjlQQOUVPb
1dH4hK4qhfgs483LZ+u8YKQOoXAqLBxUWkJwEKkVLijQuVYNj8ANxLiEPhLaeNVZq16RZUX2AOBv
an+EJBpH+zWXvA+soR/qWtp6L6xWIqh4VOgt/lvxxwDYO7cd4Q0APOSICrhtS4tZvh5z0MaH1Njg
a+AgtALSl4ZY1YvE/m7zLE9WzufYGyJxCdn8EiPHHf0cr5ExDouJTe3zmrSbFGPLJM8BVcyvXk/l
oGaYtML/pprnxh5sF4ovxPnIaztBb9S+Pepf2lDB+uxZ9zGU+K0yEX8l42VsA7vBcuo9H+bt9C2o
rWrMXi30XguUn6cwxHHrAhQ/aXC6cJixKjNQ3UIAFGB8u23uatnaIKEXWAAa4btfHrox+jlgAUcG
0r42sSuDLCAzMzaaPRmI79OlISRQLE/k6TIF4gu3K7bOFi1skERQGzWlDQx3pHucbeBpx/chjmkK
2n41op2mLbD0qGLZ5FD1xghBVTx1zqkIqWXNq3GUPATRvFifLW0UhrbI+yyyIU0FpkcDS5azYEqs
e8eeE/BzIyNpxGD6Wcbp0lIf9Y3tpAda2mEIlnfip/cSwigaKRUw5oRgcQTN1dgVR8GBlOak7XTI
vVmZo3Ky9t7QhG5pyvoEcubEbYPsiy2WORV/AI4UmMJqeC1fSC3hXGG8rvlrFJmvhbsPkbOyNpjZ
ihi/34j/OpEfv4uSE7Gflh+8uXaXHAsI3CAtev3q8Mc+vgSbcfr/LWJkqFM/OrfVBxKPT+ZxyIcI
I1wdGcu0sCMuJHQjz+ifhMazrsXerdO+ZdjgdIPqfD4CT/y/CLU0lljPEJKjcIwN5SoPClu2kAaJ
pt7KpN2+9sqBCHqFW1VB6rWJAJG1klkJlUeffilF+8em/5HxCFn5pw0wgAdneYvxFbOYE4VzYf42
fsiJdaGzR4i+EsWf1hgvQBaIl7H3BmWsHtKWI1aU5BSpA054bHucndgEInqgZP+3b5i4j0Bg9DeO
f8XuxUyRBq00+XZTgaHfN2LoegsaCKr71a06OVZkJ6LwvEyp/AhQD4ddfsqI6zuQ+AyNdm3rXESu
KToVeVdZ+f5A/gcprrnhjv6FmsmdB7Z1mflXYSOLUmxMHwOCqo2tEm/d6n+xKGQc9LwRsk3RCfKD
Sh1Ehk6BEMitfYllzMfWRVuICIyeSFhtZ02SPOBHv/WtGlmgXwK6yEJV/cGv2dmQphVzWVzl7LrT
rV7xcMJY4x4LaU3bjeBxmo3wp7GxIr/2k4vSplO8J9lU64FxvJp6kQjODjaUKe5ZgnebD7c3tJzr
0RX9U2mq18FHvCfJFc/8+s2nxkv0AcFTf6+aq6B+NYOHhJgSN0svHI3QqZCgw26ZsCrJlJt57Hm4
kTrz5J7JEVJqqAnjezbbANhPUgCCyN3i+fXFd1uqIJG8kya43eWiXHAmOWlDZ7YGD0NgqKmAzUOo
RPcrGqwwe+kZOzeKIG3x7SnJZWSN+qMMua5mMcpf9GQYK5+tvUc9rGeeGw7nqJJVbdBNPdeK/qKU
b1oesc/c4bLWCyQfsBWt3Bya2lISEgP6vZuUKetkkyemJrwExycV6RDjk8t0ivXIWhLAUA4zWIe1
VcxYohFXsFD8j/L1tEV1HwvKuKTxPlOOWl5zdAqLaR3FjVGl8X8HHxhE9uf/v0s/gh9zfxg8X53U
BWEHhsJ4YgBaW5MeCiaQoVvH+wUrtDetNLF4GoTgic0Fabx/8Pu9MdD/SYNTPsle/CqWhJ6CpjTm
zjHJkpqe4KTbx7QmSA7Nl77rlIlk3UOKUeQwHmY0nDeVuhvt5R8drepflnRyDyriYlkW+5tYCer7
ml9jzEhSBPSsDstRXKinehLRrRZbJCziw+geVv2ossUo1jFfMcXsKN3DGM2EcA8ldiN7EmEJJbAj
N0G0HOuVuAVkkBdv7QTXb2/uz/o7/msNv1n6UXq9EG25axaW1dLqyubowQekaNm2Gn7SN+Y+dtpX
dDHtcCClxdke/UCx4GZX5usfL80uAP7lPOeetjRI7vgxAprEifP+PquunoEd8HcSxnNAFlmo2u+w
qMzggwrDcumxEpGpTjWDma3kSlDAOjxAb8DnHzejwhIcrj7A6clKORsFxqyhoJuD7z02PHi2uNGM
vusQ/AjQ+fHrLUAsulh6wPaOwFT8YbqNFiEhFPXvsjmY1kog0WIifWlBC3uPOztVSG1n7iBKZeFS
f9K1MTgqpn5y1LPVWe3Tcv9H5s25sdzH+TLUujOwriSqDGJIJ2iHw2pz7oOtcM+sNSZ6TadXnhqp
ngYkw0PfcvhQiDr2VzsRqmC50EXu7GhubFBP/8wV7Veu1v3krMJHxH8X9LDLRj85qSt0eugvOm99
FJR0PoklB2yrFNLXoZf8IeoTrDpDvaBtVV+FSObFTk8xdKhvJURZ2AecOnSgotYNpkugfWu4tUDG
SXlAIwnvqvi3lYNmRDxD2uOV1EppHQqpLqIG4Csd6XVaW7mC50gAldTxHfH0yxbbCYcjNFyiq+Sw
066/Rtq5hOw42MnEOleTdtkYIDilYwqWDiZiB/faFk7X8hWQN8r9qg/U7pxLk65P00h7Yfmy29pe
NtevnQdPjKQP76IGRo7xJX9Aeds+eW9SivqRFsdW0hWogeumIcg2rhZCf6sSHHHyLohiIlosPmrG
iYxEO2FY8e5oIeupsk5GVWOARdCap84QD08zGGrADGaldntNjxHJ3n03ZplgAjxtnUKEEu1GJsK9
Vi7utILAmwDLVUQylkJnSc8B/mRLd3fh9aCBxxIjdiaYYsUjN9aDtvenT5aumpTieJ7UCl0TH1i3
+gM6IVC6Ro/2tmQytsr/5hsU5BAYXEgekpsuTojEv44Qyi6kPtYTOrKNRC9oH1PQZS9fiqslx5fx
P0y0kDujYfD9qXe7B7/GyqizE0XZnCVz9WsfvLsrfbQV6yn9fca2p9NkOkho4eCOQUyOwwaR6oFl
EK182tbz/klOXfiNzNf60aOOQY4iJj1kUXEOMCditIV6gGU3t4WqxxfaReUiBxaJm0Yj6Yx49iQT
HOWdTQqwVA4jSy8gLZV1XkHNV3d+knyIFXneAs719Om2e+o9xKCFsnE7mBckL6JtniBZqXdo4n/X
voByBpbBMPGKD0DqP1+szn/ZdRBlnVngf1CLwq6gaCu+YVDIbBNHLe220cvDy4oiIOLKV+hACcKJ
WPDWuBmGQJJcPma9J7vvmN/eKNntRiikazuZ8mLgUrpD80podl7B3ImcNru4WxpHfYuF9ZIytszw
4oBGa6z+zmU4Sy6CILm3jBQX3/Esi/DwotohoSAjhZKrCz23VVj3KddTj+xLKkL/Mzjt/M2TmD7v
dyOpbPUKVmeMJXKAE97YsBKEUddDtPOI8xAbsxp1FzL/GMSLlkwBNLVnbTlVsHzTzrY+uxrXydts
kAKWCsE9IUNuciw/1RYjeq+HMADacv/K88eraxG/eyOykZw5dCvJn7qtrDAN4dp83HzOvOdn65p6
gD+XAywwiRwkHyELAOcHjUoJbe5lX9OMGlvo1sjnkwU+1pUglHliU4twV0mxBd2k2pL0bK9nrFS5
1DIEEcj2sk+Bz1q4Zl/UaI9eLg4Sy0baRHSpNwqndMOyoW5Szu+qokUWePFINKvSJzJ730PdxMIf
a2Nr5/rlv6kcZSoxSQ9TbysgL92NJQo8fOVxyZokkFueX9kYiORwl+jtOkvFrrOyctwjS3dj//4r
7OQvpyaokc0KZ5DuANoDlz50hdjSofQq9VDPWLS2PLVMdeNBKS+wF/uF1rVdADFHBuCsHVF9Uhp/
KcFB67zAxx9NrdULSBIpbOiSTIL8OziF4rWq6XsUnQHJcdoYJzz3lCtgTqjgTrgwKA6T1oNO8KgO
clwpJoSQkbheIxIXt/sVX5NSTSy+rNszPnAAIIfSNNxwj5W/ebqY61QSinrcRyTcv+FASNaiQrho
STrzPCdZY4UfOYh2vQRWiu1CfDkRotm21UUNm/msyMa3yR5hpXHl9kg245CUbZrW/fDZAQKFdOE0
rrQZoTN5QQ8fqqODRi1e+kV6RpThOZUgC7HZXnQoUmlh+jY3PnA88pZc0mX36IgVsrCi8JtE7bWN
JeLaLG1XiMCpWGsZ6/WfCwQyzh/6yGhB8GqtNohQHiSzQigU39DjgCy7scYCLC3RlgtczSpFhOaf
/CXk4QbnJo7cEdAzV2pB805BN0InGPwkVtE735z3otkd64rw19RZ13+H6C9MReCCqAlvNRNluFO3
MVXiO5XxXEayr80yO5XhyDDv7WE/RbqNHaPL+WwhTYhMdbBoqsqK53qd+MlDZwhDv8w3KSROq6ai
wOgfuwVXjK9PqIRIMzlFzOM2oqiC/IjLK9FZm9O8jOyYAqbl1HqCxUhw1SVOUat1DBSz/oVdoR87
ccGnNQB4buuYTdjbVyC5D1RGT9CKwzOuhd+8W4I/uI+jmFNXBwrXesLfSog0OXpnpXodiHpV4qXI
2As7B0URnKBzS6ejRq/bTHw2o632e3vCFKjEqfdq3z3FgtQ+bDzFPHK+EnF5KamZqLLZ6xqN0A6V
gVvDv2X0dlk5Zgo2wxqBJ7i6vPuzU8ZF8fCeOvfXi/vyVqVrrA1QdXFHcPf6UVztY7vkggeDLiD7
F2TczS2hSQGaTEF79Dns+4c/wL856u1wBP0lqrwxjQIElr5RYWH+3fq3//w4da6Bz2DmW5HhU4a1
a7v8qlhMptTchYUehPWXE444lP8b4GbPMZucxW9Bx4ujtHS8uLz1/K4HWOgn+Z56eJMhny/q84fM
I6Ij1uKWm33AIfy0MNfFYk/3dubaxZHhrq635FWad+hfSeUWJWqLAdGcPfE+ij6//qTJy5osTDj5
oX0QGtzMSwrNz3nZGIX+Ntv9NzDJmvciNodUMzpIcy/grqajkJr9DadaZx4yZUS5UcVAOYU62ZkK
bIQCoLsbjmXSpV85Y4bVSBj7AaZ+ldCb8Vx0wkiTBUMYDrZGpCbCYBFgVLirQXnLJRvVNGpzBF92
SO7bbpRGwFh23UM7J4arpdpfAU10PDLoLpkU3Ph+IWNyjerozpjv3g8jqD8TUDlMw9AXFPXsrwn0
WbsFhWlrcQmcO3H3yITAIBCzJbM3NlfrnKtmlYjWdU3p+P1LudCuzvaRVQ0ckKlIrDXLT15royGB
gBp7ivf38BYyoZ3x34bHCY7Wd7u14g7y03TsGNQ/IDta/VaTtq6iZRg/BHRWdkO0yEy2ARJNFtrt
w6kqhUBuvLl/i+Q7nAQo78xAVNC5dkXBDdak1i/RtYEk0oKEfTMn7DdTnAn9dLpbbOUd1T6TcPNH
mAkkcMEcuSALcE06jPgctthH6teA4VXpVDnuIg/Wv/rDTHfqEvapXVidcmtTJ8L/bp1mgagnLW2Y
f/62uUMTvoVLiVEV2tZD25FfnH29yp76kGyUj0b9v/t57zyJYAWgd8JlFZKFw6QzL6uy47GuDdR9
DRSq3Dt1KOdH+jHE86da0IRtaQAG8lBynO3gDnO1iBkPWGp8M62xLmNsT9LtWSMTYRdD6WwmDkNu
nkYMC5E7DMasJG8uQM0fNfTVhxSqpV+ysiYbDX+V3ivOKJyXk/ahnF4etiwd62ATM5ARj0PBfYtV
RHKorZQBO9V00uqzCzHJ428SX4dEtm8d4awPDqrz/aryk0XMB0S80xq5jdA5v7pOYkBkO2u0DGdS
2vucmmdMsfCOI5S2CdLdLisslN6nvyxSN+H99at6ZRb/LzkgYxM/tO2r/mxJvmJT9q9zpIXEx1bd
hbCspzgSO22+touOWwFs5dbXqDAbvLV1xPNlttFfK7JHp+R6FUxc85VpU+u0KuUgLoDlS2cOKr78
HiBWqgNW8vyOUO6ISHmrokVvbIH1cPj0VBC65Tx44tvR1dX3BBkPzv8L6nA+L5OEwtCnIUVfm0Q1
4/KsViFf9EyFa1nJIFaFa6SHe5+e+2aS6k90MtNOuaEs6KuxWPiZxu4dXAuUw8K91zRhG5tUiuX/
r6ysbPsAjTPeU4KuEVpk/aJ6fBjlXLGbRIDzyZYKLpr7u9l/2c6PPDjlcPlKrC8TX16tRlvA4u/Y
rrAL6V22AAOsiNIxuBaDW7Bk8+ZBYrIYacFI3dc3r8tZlAFI8AXlL3HVlGaMyyv7SdRHueZxqHPj
9b+dpoLewggXndxCyBxUrIzO4XvLMyR8tx07CQbBZAI9mkZCfIZTloLhOdrT5szEPxVw0/qwq5YT
V7QrcLwiPQ2RlkUSI9uyKBZH4pJDxeGpVodnhTTWDt8i9V2tKrPV7r6KcndANwOmS7I5uRSkdcNT
ybiCz4DgOC3sPAbBuK+7ttPRV168l/v6P8H5KH52BRNAJn3TgfEtrYPr0zG/KUa5l77IhkuVSrCp
oGeCi57JOWZd47v2YPvvA/G+re5dy9Ury2x6TCRXo/Z1q0BI/y2x5fTnmU9EtOyvrm6Weo9y08v3
ZwCyScFXR085NOshD9hG/DL8blnGZJ6yDoH0nYW5Qt5KFSoUlZkq3pVuRb1HHTegp8KaNSrozPAA
PCfAHW+j9aRJwXZWdT0hQX48JmfyB/ZBYqGynbrpXQd9lv+BIUKWt/zxL0aFQdAV/ksKq9FDyUQV
zProJsZpP38jZC6qGL1HUMVPK1dGgWT+JSob1lh+AAYBms+PyGdtrEmc7TarpDjuvb3S9Sfk5M/w
YWc7MS9rY1mHVyuXCndXYnIjVsPFOWW4A9HbbNEMWMQnQOdV3YB/yFoQwCcXqnJlBmWOiNSKQa/Z
sKhS4pPR7wyQqyaMazdUIndV25z3X8jRsnk6J3EI8n5HO3L0YspP3JnswfRseAkXiYoGSzw2zJfc
BkCq5T0r9qJF1Fj7wjcb9wVz6ZptjxOJOj4bsDuGaS7MBVsrM3dv7I8VngXAwzwIemLGjisVsMDp
YtdwRdFnQ2+1FB3H0Z2Mo6lJRKrU4mjmY/qw//FnJC4tHNXn3HUBANezbw6VYVINBI6CsJt0tFLc
3AaDE0IFPfwyT1Xc+4Q+5fmMTPuJ2UpRwz3uK478J2HuvWReylnirWpQgIOv/S+IrBi17BT0LqGH
mCsUMJlGXUkha+WzNSk7Kx+sJ4JJfT2erwucpg9KQYL9v6hqVJD06rVfV5tTAkXTxDMx94suMqZw
cAYeHlCsIaIHfkfRVZu8ECcPUWfbT0/h0AV/g5WVXwzXDzdRy/GbEbaadTkM8+bgyadIVw4FUKzm
vOmhY1yGf84vBQr6N5/SEJzVXiedDRNMBb2/Eq72qICWona3G0K04ofPlHB/foeDv8GHrreIGfIk
xZj22Eynl5nSxxVpOR/8JQMLfQLyz9kJlAfQ/KHTDZxh3c49R/3ft8BSV9owAqss3z0Ml0zndoT/
t17bqxV2kxw9sUydwx2X2DU33W1hsDY84HYh+l0iJu645FVov+Lryhcatc5H62COaPHSqxHyA4c6
DhHsmsFm9Joj6rtlghvhOyTDZUb2uAbkBvycyu9adzfPo3P27R00oCCrYBnjZcBoodxT2eXW7r8X
BBKWHSE+q6c8Uk9M+cZBATC+IcbagICN1zSjEce8iExl/uPudhmVJU5fFAtfxacXu59kvmKcGymj
KwOgbHfBf+UJOaj7/Fv3PysaiCC4kSieb/q+iad5RvxZCp4y627Mc0a6E3eEfniwkM5A66PZA8Sw
Kn/41uqa3wzEwCBJO6y43KZDN1nF689ErI4YyqpcLekI2XPQGx4I8giCsY2BXbYo8dnM7Hei2BkT
EWmHLcwjI8gTBt0RZY0P5Ihhlxn2yX7OV3dJHx+rUjN44Q1lG2po7nX0kVjGKKqjWurp0ddbD1zg
dybPRTAcSqqwpS4/vf3GlG6EwmP1Tt7T67+AcujDBWaV5xPOoiocftIRszTpGespBGDsszsUK+nu
wVDWVpmTMMH6CBNIewtR32dntgOlH9DvDEOA4BpJzkXOiejsS6Ki996G8gur/6DQOygRLIg0opdz
jMK0gr5YWdaYyQHNpPygf0+/U4aRXwHxcGQMLO6uK/pd2CaYCfz+rE4CoSWSWuwAXHm1GcTFfoE5
msYHVL2AYwCcjRed/XZRM4SwUxBkRuSB2689lhBAQbyX03M8TRlWgq3ea3gmB3hN2zLYTGXJRRvl
ZFvbxiFR2jWr1b5W2Ji9pRrD6ViFC9pjJUv7XOWJHbh5aFNkE9yP3pP+Z8mGlaMlVN4yKLLbS8kh
+CJdcpKsmiUYWJAHOy314+7Dr0+m4de1M69xEYUziEawQ3pUM8HyeymnNqjTqQ0Ej+fUc8pnF4QB
CEHmSKxoK/gD7TZie0nojQpnh4/5FpKthWwiEcxBPFu+tog6Nkiql+lUBS/yWDGMLnA1QN+N7GaW
fYue+nXUC2rW+5L6DELRDR/bAnKS2CjwhwR3g+AS9cMd8Jj+nO7VrDcb61UXNeMFLpOP+qBg60Xu
toTnSBZCfR14ehcSTGNZuGALwGubkanB6WJ8vG3W5OoyLZheKgSR7+aMjcE/hka9oLJbuQNTXJAO
zpf8IboJLQ4rx8E7kpQWb3A2Ijib68MdkxHwQZDIDgM6rekYO085CqqfFrhiuBqOTac8Q9seB/B7
vNnAAg2mhngTvK54OnC8XCMTTrefVKW22CwcasNeHn4poKFAc8pnR9oFTIoOlEuMK2CJyC/V4h78
MQ0W6n0ccXVCyhkq3vGBuRwCvMB7irVwI2nLur+YD3ZmaACEB38UN5bqpgjtWC+aLWAKu1rn5H8v
TLZQ9g0C9spOV39wYsVqCbkzpk5LBC/V+X7ttOBE9E1Rw0dy/9q52si4NzkpyjrZGhm4XziXNdX2
C++cews4Aj7MMZh7NSkgTbg7c1CEjl1uxwO1c6QJ44hJIShKqmy/li6UT2CehqJzKn6t4EX0nNed
xoxQRnLjHkdPBusJEDP3d3lXgFwN/jBlxJFKrhRJvIwkPHTWGPtmclbTn0DuBJxO2DaL26LYiLJw
rzKWDpNF4zxITcCp3mmFc68Zh/EkpTo4c5LwRWm8GagTxkqtKXytHLtgqLUaMpzfw3js9hfCSQyX
8XLSM+aUkm5b1i6qRbKX1rYtkcRGhJCOqgu8xqahhfcb9JpSf2h7ENPSJ7muEqt1ZPdyS/iCuM4r
L0+3+PsezvQwhlZyjuLRhFNcFh4bmxQ6F4PHUjk5KWZslbQlPEirSRUCFRmkWfbRF3g/TvLIxI0u
DeN2ne+xOh/cPaRuNG+032N2X2h/bXzihXWr5Qx2V82nUq/X39x3iwtQuICCgeO+YPrGzJhG5tlk
t84A4S4sXemx4oZjyA8xA5k9UNpB9D7HirFKL3iD4xKTVh2Z9QDE4xRuT+28Va792uzA/rkPJIbf
qpSRQdVD7zYyOEOaWlC6r5TEF34Mq2/IoGX8r/5Yu4N8Iv6Sm+U9c0g3ag2kAAsYLw9xtpJvTEEA
l6CAHsmh6cZMjRD7TBTltvlS5/deJGkFuUAcSSFudAj+c9HDSQi6CQb60JfHvLG465T+ejqtepCM
R6J6+rGFtJ63KXwygXgyXPYOwGYq2QbpvS7NJPlon9MNxa2JzSeKKeRys3c9ERbPDDGWkPHKebEZ
AsNlwuRcaBdXU6xX9S4b3qCV3wDm8EYLpfVgnrdt6FSbl11bzoroz10n+LTqfgDZBnLAzLuWPK4v
JkwNcWeBitWcQYB14UK/Bwt1ZJRmLvCkylKvBvuyY2GH3ODLy3ZkuMZ03udEUmP059nNz1x/fz0z
xo6n0yP7lY6trwGl7EKAqU9bye8w0/Dl4T0sCcS3T5LGOIojURJfRC7HlmA88VS+nckJRAfKOAwS
RVIzLNwEelhkP8HXZ4IZa6mjJUxw8C637lw8lyrIS9wQXyQpbRAwtO3LWkRoqhqaAiINNzAKxPDQ
g5vwlRhFlAzimRvaXVYJLo5Z9KiBfLvJnb5Uy/HNx+GAB80u+pIig9s3mHGqzAFdZiwkqcsXvGsp
HP2RMHnD2Yq0v7DPrXwVtsYtu5iCTnf5apbOLBSPutuypHHxtGdhHkvmKtu8Rg+LwbHg9E/RNTlm
vt/4YLPMli1xGXUkMPg5rmBJfncVp5F91jB5fHdk9eR7DlRc0JRzqfsgtn+pehzH6772G2aitQn6
K8ux76mI4CmojQtUoF473iaIKwQMa+XOZwCFYoq0NzQF9maDaviNNwaeSgWknm6oe6uZ+7dw9FlO
byhtMKSsy4LImX01kDHRxdB/5NXr7Tl2e24RHoxb0EIuxaxFXjADSBhtYNfePsYMbpEv/4UroBHu
YRrpSmV2akzH6FIAISxF/KVuiWHGPhoMm94O+Ti/FcW4jHiNj7+SrxYB4ZU3iO4O5DlYY5vkZQvW
RmBC7BKalpWMeHcgQVuLRbTQdAtGjgGrDD4cKwSoap8Zh6Tf6FdWH+M5B5GnSaQsipUV+lELFXq1
BOG3ffJVGWWM1MiQXTmvdzeZH4Jlx+B3GeRNvHnsS9X9WVAdHK+JHKRFoD4v0FEspchpQlrL0Aj5
a3nwZgVdbLsO3T6VkzAHCtL6A3ymkbCZy2bsycu2yPJ1nO50+3Tci7cWPhFt+bKDcvuSqWdKu8a2
op8iTfXfuOWSL5l2yL/YuA4gV9+iNzZDClzBYuw0jBRbqpdqMfdep1TrIOXT7/4wGabCgQOTV5FY
vAq/2MUNiRE5Lg7A2nQietfgP/D4PNL88u633wi09cP7W6VaDXfwfmhzCPwrykUDDYPhpRZklras
xtsMY10w9OQuaPYtVbHdGFUGrxg+p0olh/J0dAFMU/GTRaXEnVV6onxGFibl1JitNBFS+9+jKDYK
y5TmMZsB2yE1ZvGxAL/Tu7XF3n/UHAvxHQSO/h3f2g3SriMcQsiE2AaL1Dt5YwWgsdGKRVeYlAl5
lA3ouLT55XeFV5RO1m9OczNsaWPECsxUV1z79F7ioDHZbl1lTbJyWHSr1UXHAG2Y/0i6bX7K3kg7
sgBr9FgvE5iYoq2v61WoSsmodGKFfO9SMFpY8L86UK0NkvKsHlJzo1JtzeIrUT61y4DB57Gv+XUZ
tcu4nqv+2haCXAuFdS/Aceyo6FQq5KijaDNeQ9qbCAnOSuWHxsLbYCmJX0hsHQrKh2ScU1jzL5NV
4oVnEin9Z+qpmMk5YaGCezB1JC0mhX58kEiBOj9JAXMly3HmOoGZI8wFP8bHp1NuJc7+60vnESZC
ghCkQoaHxiCEpnDTO3Hc4GtTGbWtbMlZSvQSHaeCfjC50auaeN3IuGM0Hz1TiEcWEnGToOwXPWyO
i5Rg8BE1sb3A0Kjvq0dlUf7vYO2oKEtIDZO4UUKQXSyy9k4XbodAZg88hRXs+0wnLizjW0Ldjwrh
OIgsTqEln/KOi+xjhR9YEWBZ6AhKAmBgpUMmyD/9gcUh5xUfoIk58ImklC0QAKbJhr923DVGOH6A
WG2aBGfq0Y9QIPnqtZ3Hb81wjktFBAJGQxiXHs2YlxNhd4gNfue2UEzRLlt3rjYgIl0B4UZ5pybP
DflI+QwEvCspzO5SYPI2MzwMuUj962ol3Z/szAQ7/e6vv3vlUs/4V0JCwtQOpHVrF0ba7PSw12Yd
ZHcGJC1lyKHHGllW9pnAxcuIOnREOymdnycYPSWiPMzxd2Vq9oxr53Cd4//7DL2SaiCQ7cwKKeH0
SOJSRicdiwiE1Y9VzN5UNdvJ5+n8TKYUFAIxfYahit8qiZA3jlwS6nE1fybJtbREpxvRO4ny+Avw
rpJjy84/lsQ9UgXJSTp6S5n1lXAe+Q5zDJq6ODkLoyCNVT2+ohOHj3I1pdKvU0zJJ4+yManLldFY
mDAPFn0avNYrDIH+1IA85t+H+MJOVgeZanLKZ5/jXowCVDfblBWjdbwKfd37cYtlHJiGKfXGtdJ+
q6fgr+PlrLe+ZM+GnbixVfxTIvOq5JFqMz/jRdGtRqQQUsOnVtpSOZzQot3WfnVWdbZX64WUbers
u2AEF9IC6xtiE3St4FH+t46U4o3dRZtj6ElrnR6NgIPDQIHug9JOSlgcJInP4SsaWBDgh13/fOoQ
u3A4E1cljyUficmjhwJbXTI0HsPgJV3UKdV2oXkZCbxyCHM8ipUde2Ju/vIM+eu5oFn7FflS2QHD
83Cxjo/i8Q0bsTmnjwczXud8lLFfRBrmGH4pW2BP2zORPUzoiuImeBT2bghsi+XO5DydbsJiSblG
7s9ydcHpsMndXRhTu7vPdXIsrvIQOUsAQ9fxP1ZfrS1vNNa240aC8OH1Zu+z0ZptxudO/hCaeJAm
kWx2GzC1rstNmRX1ND4DU9c2JRMwR6DxKitEuT15ibs09CuGreD2jHOxn45qPC0JY6I88nPvlslV
D4rC0pHza5gEbkrNtjNyeZaXztNd4+IiLMESCIdxWjNrGnVrvDeKff+1lcWYuKuMNWXZsBdR0rmY
6jZtIcnvBPACc96FXxlVp//U68Sp2sxTa+dbIR6q6ZxKJ0OLtU5mAsMWIY7GJiEO7v+XU8GmWoD7
wX6UNhcO3pSTM6YjFYCaYOj8c/zPuGQ6efIVuyLqPs9CpbutN+efgYbuvCu+RC0/QAnsabUj5v2O
gxCUiafnXYlq/6ejcTvnfypoPDTNc0LsqDRzWnxjQyBo/TY7mTuMC77hsNtYPxVE9Wbz3t9mDAvY
+EadnXQDLXfFZT5DO96SU2GojtWBCjdANpHFyoIowgD+AvemIKfM/rEuCpl+AihE1Y+GoUUDlOJw
vQPYc4KUjYOy/mRZ5Bv0By7YvdxwJJ0wx2r6+W3+5311OK0/0w8Hh+x/cbydJ4AwnDPWFh5t/mj8
Kb2M+t2m6qINz5YeIUp5v6RY7UIt4f2YHFHmfgXMT7eDXhkW7kMWgOqCclQ+WzhHpLDIYb+nQcJ8
VPFJbWsMiBQkXdrI8gTJssVdtdNWGjCHMabi8IbQyVDYZPMFHa9/SVceKA0JitxZ7mYRZdjsy9pQ
T5lsKGcEubNgSdG/GW6xZ31sSTVaQDeHY2o0dV/KUT02/O6NKinGXew7DSqYm46ndHFoiiIfHzCw
ii5UFtp8CtijMBIs0UZCPpM1RVdHGqcQTFsJb6FufjeqBdPcqHKutD/nWFPX0cyLqgokDwK7d62c
X4TYla0JvW6GvnW5xj2P+WwoZM7YhL6yfja/jlOfPQHKfCaAd8hXbi8DpaFbA4V2mCXMusqbyJoQ
M9IqS1RQ84S6HzASn3CDHaiMpPcQTkTzWvsaLjvxShHZrJAbtLKwOUvSPMoW/51C+jB3Miq8NxZ4
WTQs52nqZKZSkHkNVyKo9bNSvj6uKOyE97N9+z3aBCRmPrOSFrG1cXhK+XxTSgZrjD/lJ9GY7E4k
BKmbHIStpeGcc6b2yjPJpDTXjERWqrQeFr8a1dojgbOB0Z/vc6yPFMLh2DbLhXJoY1MJreWLtCBt
uULNUxz6AenmSWuIaOvSYOVCEeIRXYMhbEDJAUsvlS3Zg65LZDOtgh1xzTv/hNrj7NBCyCs4Tg9+
+m8PWWLAW23kxvEJbjWl6XiBQPy28SjQ4cuYOSpGpFPXy8o2ce2lydBviwRnh8HiJ5RvcowtNypx
Edh8mpaRAWHqP90X1nHEiFdwzZ/Hkw0KM4QgveiI/+rNh7mvdvtDgwaFPIopFvJ7+2nNHVFrgsZv
sP5YZMXlfxy4NRZKlvJwunQVGf738oH3iPcEWauPjj5vgzTBnj6pkDXQwJ67pD+fYYHC92mWQZVa
xuUUbBCHVg8ok+VWPipL5mm5UlFvlm0X4MNxqLrL2xMoFXt1hfFPLrJ2LYygDov0Egskj0LIWf3O
td+zN1FbrxAZBeJ0LXobd7i3Cyu1n+BEHmgQJSsZYja76GGyNgRwHYwAfohjOGPSqYz8CXox+YtA
glZMO1MOoIhbWhHcV9Tu8A2J7K2MOcuM63hef2K9sTsjmCrNi98Zj4Ji2zHhuBXFOaNoRB8YJ4em
Wh5T/+3B5zShBB4nfHIGHt3uWT2mo1e8v7NgckkkmUpIdDV63tHvGLohsAydNLYknOH/Zh0NEk7b
IZEkttYVlvlcfKXPiCkETf7YiqaL2LNEvwKS7X/U/MQaEI5dKrrpElxIxPJhM4omUpaijO0NIhQQ
+e92CfrMkbuDAkP/JVWIi/ocAIgMyHXixjYUACHQazGhk0sJouh27jwo0Ahnj/9H28umerI35lw9
sKEU0oTkd/HIyZmPp89eFeCMlHstEUYly8jIcqibWj6fJpBgXDdPt0HP5W6E2UoVzfilhO6cn6S0
N2NHJk39K8EdXT10nl2XmMpN30tb94z3fSrdQStrLVfogTkQlH3s9AD1ddCrLgz8B+9BAzgV91BJ
1ZhbxuOjQzDo0x+kXJr9u0CAvtSV7D4l7xWnJmBvkyS0T1oAp2OoChh7ajlayLiKHkoXfLn2MzAJ
uVhxPxxmu+E5ewn4PKcZkQPupt1AjhwkaSnkIk7MYASgdYd79HSp25IIR6Q/yX9U6vqng7HPHPBM
kxeuk97iT4sC6pEIkY8Ogoq7y9BsHzGvofGpr4su/41Sf8dnJq+lx0GtL2GE0hCukfRwNQYtIgap
MVEjXolRefslK4Tin2aw4IZDppwP70i84sAK+Xd82teRi/b0ZZ1bJVV28ZVT5iOWa1mwrxUklg8U
P9vg7PLm12rD6w9ORD7hhYtUsxaRSuMRbeaWgUX9pTzsztFDN7QeVLen46bTEg5kFVoqdYNjy9sp
beFrjBJUIRUvOP9hlapt4+YFiRnMTsM3wzQjD0xtnVzAddQ/CUB3xdOY7/kpaHOmL3okRkzjnd3X
k7qocwhnB8NdFADijMos27BBtVTfvEb72EX3h8kPXUDrHZO1xP9w71k58hfyoGoKlkdSSZJw/3xe
ZmV7C15uKgLFcs2drgQl2jnYcpcFuw5HaC3E+rjBCgoNrX8fM/g+Sc3TVXzEHqaHLNryIaqruG9p
cQGFO72gTCnLwBYx6X/ZXWNVnbONkmENdu2O4BWUtu3VaNt7u7cMIoHbZVBMK4o0OatsidIRHlT9
0igyT1sm+XZ6JK8VK0XKZ1uZLmviOX/130fZD00yG439Nw+844bYbFgpCKvmzNLIyXRV0ufdLiPj
Ek1kcmySgQab/EqEZvJqbSc7NKXbv/XFJixIYrmG6tS0PxBRIb1PBTL1Xulrp7e02XhlBt98Zin1
eRq+4JDBQ7myWAHdHFqyoRBcLaZ1FmH5OWoNlKLwnR909TCuNON9P7c88Nf1rcvvITMVsoUaB7Gx
1BxqSRkO9ox4mXUClzn6oY5JutC4tWDlteyyFkdfr0TsWTkChRCZ+XFmGUZ0FiwaPwI5+Vl1LTut
hKiQ+ifnvBW11rVV4NOFyDxl+IDyWroEz4xDO+yL/slss7viF/Dm9DMBjjUQON+J1qWHxkpnzRO0
6J5dXvSNAmWK0uv0XnhUBrMqxe5KfbvUTkkjJtA+gMARP4814d8I7sZD3RaVFf4YkuoWlUnNOTaN
ZOx+9O4DHd2q9VgDXeCgk8gaOxn2kwu6B7rUGpIilq5QYc8ejvyp7L0xeuX6fX9IpBRWhj6daXIR
WPuCsFLxwC2ahYZG5sgUH7w9Vi6xNeP8RsdQd2fK2B/4q+mWeBtTFD+qKEuYZNAdOt54l3eQCQzs
QBr26CeBQW6Zu1VJkehZ1XoSk4kZhvLMxjdT+b3tKFipkM7hDrFbchMUuQrYQIw1oESe4IAFFvx8
SqQWH5br8xfSWW3dAv5KDonM0wtZ2k5CI4mOLC15SMIPnuNXkh5TCK/qd1iCM9dC5aGoy7dtbhJt
3FfEFon1JCJjjCXgEBVlxRjn+Nwo/+A7JQVc9F3GIVIuaZKeWcP+VKvK8dC4YypIXqPeTIjPNNWu
JtkruWhEYMz3RAJ0/ipbXDF0zu/pAR7CZ4h5OKOh4LBJoSg50oXwXXy8w8JV7nXXzaHl6rjmF7LC
HKCvdThiTtLrwH70UjSDQW3xkRR/eIsDBEmqyKpqgO1ZGx+6KKYiK4o4lp5BMEibTbolUl/HHomL
bYDR5UUH5g+Luho2Lm4EL5S58Pwf9jvhEkTfzTda3WPUOhj+54yQLGeQBUf8JxFsjNwjUnRuEPbb
8V4tAf46zfE+Nbec+n34Z3VgsgFghWq+Jcc/IRe3aOHOtXpgPPQ1L3nHmH8cWGXF7y7lIdGXKkHK
KYwGY685lvWQrF+WPpeEkDAzbx7BmxX6CHJ64ush/HRLTvIb02O7Zcsho0bRLM8QS6QbBafBERds
L3PHAshqxAuY3q+lvZnc76o3++uz42DiTqodpUsBmTy/Fc/XZPNmufDJufoY/rNQ8Q7jOr4eeXro
RTeSJMLNIk+xlDROtKcSPS+J3MDOE2atBrpyHcpPjqOsB1/lRwk1cd3NzO+i28wf7l6AgkQjpOJ8
0VSov3KxF8CDSy4bYlbsmcQflc9JxfPc+1ls9aBfJL/boTAPyxc/zOrB7c0jA8qdncno9OVKUWRg
Mwdjt5p/SHh9Bz5AphC3BmZiNOrwkh65/l5IvNAAYW5ls7htshgBSB6yBsc9oRQyu2nVeAEDxtlN
h45/1bs2+w+JXz/qTgIlswQEGwtIZP0s9rzPkKdtdSLiBH9yvkJkBYGUP2lOR2RnZTuFpHMXJhC2
jzrnmx1gx1fC8EIgms00O0CAMx9SFINGLGLcZZrJqks8O+m3E+LRcUR82foftE0J7q4UgX3jzrCB
Wtyp5ExHJmcYOA2KGnXU76SLJLAnRENXJWmGbGmEl/Fhruv9lcDfaEQhsxC615I7p4NcAOmF9mG1
MNyCUYyEV7EmVh4fdfj3c8rmRzFxnxwBKxTHTWbIL/BT4/qTrVv0XZwqOWyCyRnrBaR3Zjd1NF3X
KR054bl/ED63v3dCy03IWz5toxTFJZuLPhKGJqGZHAhrfQByEXv6d9xCwlIoYs3ckqTGAq09Dmqd
6MHJHzFKZVDF0EZZ4x6CrbOMs767bUbTlcaTKFH1CruneQFLr6C134asDUPcmyeGFSK6+LDe2qJ9
qHbdbZ8MlkDZwP76zfHGZeDX3WaNUXrUf4bvCsV3JqJidJUOtwGl90vGyKIYr0dg849w+IZrrVEY
Nku18yaZzi5oKURBVZmyA1eUAWzdDu0dkx2Pt36xnxgp4qf7jERagriiL3o/4azEk/C66p2XzSMw
+MVgbP27E31scdQk0/eqPBF+70ZL9jCU3FFIxlGIdw0VVBCBKMeaw7l0s9y5pcBO1+bTRN7Bgg1J
IbjDNLZw7wkQ+jY+SHLnWCROQCHdiCQgKpFDTxjgnnBaCQHZxp82YYY96a/BpZ+l2vAxuVJrNF8j
r/Zq0sfjD++gwAW/BXX7gMNgTFz6d9Xs7TWjf5LIMsTZlmbt56rGhjXsaborgAUBCdfwW9pFd5ZP
/dYHr+yXW18fEkllpTQJx0fyPomVs5+1TUVdvgDv7RNkKV8vrZ+MWfW6juFaW0nFXviLRZSiVtfa
HbRpik1ZZ3oASdPf2pl5Tvkux/z2BbOMN6XPiLqMP8/9Fxw+5zeBonMdb1U9d8pJvHx+HiFGzR1Q
A1JTw3jthiW8zJCHVVpLxfZJKgk/4eCJItaDCzgW9S8S0JqlPtwAsq+a5GjCKlq1WI4TMTduYaCM
5whf2Wypof0PbBt2069q3zFVafG16luQ/dF2Z1NkOM4RuaRugKs2uIT2wtVyFhMwE8wj6F9ftsus
rAEQqJizBCyxN189SCocbUJtz4L7TG5fimwxb9vWOGO1iCEAOT/tvf8VIlnmbTtoXhSUqjl8ueC/
WALTkN/tqNnu3rwXtyWP7VaDp1G3y6nY4auJy6114uvncfCVmujjXZ1UsWTe1dEKpEZji78AgdaV
jlgOoF+oQFhgwQ8EV/KVbtuxS737Pllp2onkrS4tXmAllPUjJ9EfnOOE45PE3hj6TyBRPEwBS99B
IW6FjLr3plmEJTp21bS1aazDuLJQBDURn5/qswtQ/BKXAV3tTr5rLhSdNgQDGFQatlSyDmgha6/v
ZXoWkTcXCCMtTkodfkiJohr0UTQPcHl+N9j8HUj2tjoxAcdAehf3BcHRRtusWitcYx8jcSXI8FTX
myuwGTkD/TyQQJC5yC0CTeDYF6xbgArDosjvw34dAUB0d7+2UBlBqbS3XjcgmUP7g7eVNE+dLxs4
cZibZDG7IA/uSnicnsCAjWJ+ToOxt71wyA0zD1PDAzeB0UrITdy0Ma747IW5/SCv45OjvjCR6M2E
iko7qGD6fN6G4Vef19SPqtjAExzt4VweNOMLtPPbj9urYBVQz0DJH7ZUBMyhlaMlSTGS1B/ub5ug
jlcFY5FwAlndIhfyHJ2RjyrwBXSxFfsaTJOYCc5euzwiygo+OsGOuuVwrDh0UUcOFnq8gw2s+ZhX
k24peItBas30iX/8ATosO0Kl3HLRbjFqmKDoU5RamPjNjhNQPkHOkasdI/F5TI08UfQIyayzCEgq
bIFGsyCvBPyOSPD55LLj4Npp4kY0MMm8ms79HWu5f2VCI4DrV3J8/T/7B9mAWIfPrBB/oqrRGmo7
3UGkVMUPHbCaTdAIVYvfZudi30fucRD+o64J91agO6wjZxEfiIUWW4XmBp+EfSvvgHiK62vOMSYN
+C4f986rAXhY+WPBYrQEFiK8XweT9p7r2EptDycCGc1Dhx4F64vFZlxgubyi7brUXBBeVRAqIJfz
Q+cS9fO6ShInISYNkAfuwLp0tC9XJZPH0rzLlQozj12Hde0SJlZoenWqWHDaeHrpjumQBsCCQibm
UxVmmMzEsTLDoYCk/jYKFDeQtt4l+YIqs/L1p419TxnCUXMUjNMSlYwK8HRpCfNbguPxSBIT06Nn
lY8llFpoUTez6K27h4bmUDI0L+JG3t7H6cUg88jq5+3gvE8C9SHdy5p4SIPINVG7BHrS7Sb7UBfV
2fVd0wPzkhB6ZSc5cerEnwgGyi0XKa4OiGpoYk69BunStNmLTYCcp8iW7nEU0cA1SnhoAic2NRJR
BAERsRA+xGI+RKGlU0CJ3vpcLDIawFGy4LoxPeJ9h8XhPDnC0tJQF2JoiYlrbkKDnnwS36t19FCw
Hnp7vJQuuwuBWPZELSwmVQqNna5fMibSPRroyedRBBwKcDIlN0bLORbEFojTCZnmsjp1qdsVqMPw
fPPQ+uJP8QKzTinARE4jdw3yhgAzn3FQmY0aFvfebqR/TiFR6YRMkPMuk3eZI9et/fT8C48hUJTQ
Xm9zXEMQIOG1lCqG5RVuWDWj0xBQn9EnbQ9Ty26KEsCRd5VWPLOkVMdT6djKffcj/tEZZi9unQZO
uOjy5iRb3jrF03tejs1/XJgHTaj8iaL4FEFJmQO292xctwrOO4L2e/ZSctNntQ4TkPwwjPrmfSL7
qgM2vMNFTlJwLlBa18JRat6QI5OeJr8F1L9F0ar3YIP1Lopf9iKfIPqK2LanoA1N8xTvwDgjGWN0
/XSEzzwHZ4UPckCQOiDs+kwFFLgVoYYtQkxYGNEXQFgNCdgVC7SISBR0DoD8N+78XNSZWhKSn2y8
Eu37f9OXKaFp3G4j2cuS6WlLxY0wNF8iJxr6uAAXSYXL0VNXdspyFD99O3Fphfu+LymZRAqYuzKl
Bd+GU+mco++U5YJlFnjos7Zse64TMfwo9DEv7tBEu3OdRj65fiTTW2jkBbG40893EwjywBUw8okg
E0J81lFSXgmx4ZGMkMzfMJ+QMuoLqD7rrZubjkT58CoiCsrlXHFG9JVxFUsQhEPIM9NdRotxJAzO
tBiLV3eN9pvjhHocLMEAtawQ8HGJClpawxSqmI7o11eYi4GRvAQk2kCOjoRR/uQ6Dt9AHQMO0xav
2+0Xv6G41F31AUQttvF4AKGZzx4SpRebdCQLlw+zDcsJtuWqkpMiCDge5xJqalJkrVBU8PCk3+yx
XJeePGSIf0UWTW8s1IkrL6FJe2ttnei52nQiHyAB2BORlvaNOIA3ClU9kuYN5/l2Ow8/T/eo+cAL
YZghvGKkLeWdvmeZaic4oHoEYu36ZL7gMYAfeBvf4CKkY8Zl1uzcF5S192bPWl6HVY9w0mOPMMor
nNfAEISemngLLPorT6jP4toYas6NT0Scxn/g72R7+HkYyHCnX/ZECl+9ckUIG7FAdKfXFQnZRdz9
DogRrD3v8GVVIbv2rb9Kt2xkKzyDHXzJLKxIw7Mn5W2CMzk54XPHv7sViN51uHBI6BLzulUA9S29
ifZ9L4TNmFf5GlMT5BuJxd6hhfFhseepWrOP0J/vckXAIJSVOiyCTwefZqkx0tf3g2qzRtaQksiI
SV+qvt2Hdq310g8+oHvN5PfXW4zIVn11BHGav6VnLeyq8Wq3vHApXAAX4mjNXlFmucHi+XnDo03k
b7Fnh7XvVCXIN/6D19jwbJFW1JxMVzFGiOtlM96m/IzbWPgZePM7xcM3Y/q0K7O7MzaGcJdD1OZS
8ZTSEzxy8GCJUBfMpJCnHDIW8qsfvl8mbNZ7E38P4ErkSHDNjIWjKxisuEKMjWOhl46r4Bxf6x5T
hNsSu0elr8WwC6JrQHhx8liyhniSbNiavQzse/sfwAXSw3y7rHfFKjOoiriMIJqIz/Mxya2hKAeA
Yg46VWu2gnx4HWdxUo6vY/cTEa3JaPsQhBJCorbxNHrk0//ROJRlxc2YY59vE6jUFmqP+S8FbP+z
PGPGqfWtJU2li7gapzRp2L/iTtiLtPIeJfw8dfICLLcSXO0+2Eg3zJN5grMcyX+Lr4dpgtkVZHLh
jMCrMWGvBDDSnxMypJPdfsGNnAW941kg0a6wnojZTRJ5GOL7Dha5HntI/JdXlrZLWSrc2YT6kkn1
5ZpyI26tlFcN3YRstiYwhG/bxPVu9gCXRx+nUGl6GYOa2ZktecaBvR5ZNivykLSp6uOQDbgXsEZ1
6VjdAwwSe1KP5zeW2twgCF9tN/sFdHeCgUvvvmrs1I7FVCZ1fkWTfngtPuBIezcLoSg2SDBSwHpP
DuJwAMUx8lqWw9AVQe+iTrflpyGetNidfrmeaGmz+2T39AMg2MoASsmhMeofdOG6GAz6VgmP0JLe
8hBUA7MGNPGyrTTVnxComIixFLPVmG7P432s7lcBKUzQc15lwBGr7ZLhPjulkVsFEzKLZ3+azpiJ
dbo+xle+f34kC/+fV5gQ5UyPRAWBjJL+lpwYy+tYN/O0MVhdZwyLN8149/ayr8Hk1CoYce0evntG
TSoAS7oJ4cv0FeMJ9qw7LVnG7hjTHmS26g7Lny8sFM9RL8vhdiEnRoAgoxy+0nbhPy6QYzWBJbw0
dTwrTwvfJ43oBaTSGzByj9z8hDJSIPsHdobhj7X9NvvZrgvUEAGqRNqMMrGXvQUK9ZDqY8kD/r9A
isHDuR6w5O+klocB3f3OzL6gZPL6/wOgK6W3IhoO+aXSLPcN6brfYSWmzfqY6Submj0+55QIByEW
oVYsdsgV2/tllRf/h/IEFhBHeUwVEVUZ0XVMVKgpYLPmy81p6fAwvxGuBQz+YeYa6kJfEQ4L0fF2
3zTn8wzW7/FmdMAibvNrLs/3V+Ms4PTQ7YflLAw6dHT7JK7Af5/04Fo7NYMI2f2mlZQ96yZWs7FB
MwheTThOhs4q203P/9rfgTEfvzYZAZsv+6I80IXl4MuP8xYSyC+Bo9zGbEqVLPtMej8MkXH4JJXu
GXs1qj8C6Kv+q0zz5FhCC/cA6/BP33GrB4gzJVZgJ8rw8unEOm9bUEXINcMvyTgF0vJskyGeMjdy
nSirA+wxkj6q61ffGCkc2UAlckJY1KH0ltXsLmx04pAYfIdYUcPzgaaIaC7tmjWNmMIVu38T+mrq
qvjBhBmIAiVlkiyXRR5w0ghed8gG8MoUE9qiDzNBsOfwIid2SiGkAAiqYunLZeIxrjoixiLB8lOc
yQ9qKcE4aERLqAkodqJSJQIU6hbKgHZbA6XVqKd9qbxzcqc2OS79ETqucHDWZyiJxfUDzgFheBfs
svGl47C1QGMp1OErKlLr54NKJTIRoR5h5rBdw/RnDRQrT6E583vFJUVW7LQ2vym7UxnB5JlC0wTP
QesbP7YmTtN01kGm8t/5prz2/NC3+/MJkg4diNJw7EWs958qKWiMQ/atgB4YMNl/33q4MDrT+5qN
AxW6i9E8EVA1nSrt50J8ALrMJYViBGSyu7RsaPty82Or3+gBcVpaewRqQq3/gKBbES9hAPQLXh0v
j9nFuzV5FhFzJ5dzAPocPEItkolUJGsYMxXoJ2r9LEDge4qSajAELMYiunJG059OEBc8dpnKCBwO
bkagsW3BEFcxNhtI5IXMHfFITneob1NoFjLTrJSU9qZV/8+FS1o9koqGHqy0mZF9FvoDj2umuVyz
ksVcrpyugAzOn5MF9VykjWStGuxbMy+O/1Ehm4/1Qx6essMDe74Rs/uuW3MkmfuC4a5GLfbONpoJ
RCxehY0WgDFGJGCzhikVXIw/8EWFgEPghHNru3ftckcQZi9TBJuMmhH19DzEL5qsYyB0NaAmZuTI
K5c9IqjcnByuSaS3IHMKwt39nNHeehMX82zrSvOrYrCnDXVdAJuDp5dNyXVK/SQZTis08E524LEC
w6XwTsxmj+wYfTdC8DCvojJbY8RsGVXFRczUkhlXA7/NI1otcuHqgXGtJ/uvOHGZ9OwBnVFICl1a
ce7zg4kF6SXk22aJmTCN/50GOwJUmg0EbWqDOgtNz7j39uiWdw97ziyfFzPF6Wbu3xHvvRPPFeYG
wKttpoyvEdOvN9BW77QQVX8eayJlB0dZjonIPx19bvDUIcAzpmENyA5/hedSv1/I6Q0RPeiroaOU
IK/pkYUTncqEbL2T1AvUEGzObWYXSO0/vChJ8PG+byqWA81qWCupXwKxepx22zmCE9sXE9Rbds/n
WvwpYb4NsQt9pWYfkvttf6HdbPXbaO/GmrdJHlqmDcRnTiQUE6e9AsEEru4Y8pGHcQoIBaFCArU+
PiwEuMywoZQB7tsnCcP8HtDjgx/TtkU1MD8BlIyO1olZpIs9M25CCg1cj19+zHNIeEYQTo1T84p2
yr+vEbsyKpGUUf7g6tZoxtMuyEvse45/7doC4g3SUBcCt2SIPlPxq8cPr1oQ+xUVFP07ZwI9m2LY
QNsYo+twWcolxTQqiW+5sB8ddkytu6jXMNbLnu9CpBC/llkKKxym5FE2WLGpJgZYODXY5+NAe17o
fbKVNtXNZHhLDSB8L0dKiB9mPPhaQwcWyXbKwCE9VLPT8KggB9r2iWDu6l5CBQSXRZhhSTe21s/P
cy6PWMi8xO7NI36Kg3rXR/1lPDDMiq5csWkgmrWd0sRugZ2eDTZKyCf8Zeh+5GSUHJ9AGbdM+A06
XhmHoJAMBBAI89duoFg6F38A17qf4INZiNhbffqngcnqfF3AsfWX1S5ZAVe2dkrXpUGrPn7b5XCp
cFzFqHfW59YlBP0SGoDyX5wLG2ZRwdhZMfeXXrxsKKhHp9V+PiL9VtO+nE2n++v8OOxjPnvOt/eq
WauJelcPtCsz5ILlFLUZGP8I7k91vj4uOKFHeHyVzTRjnXopYk9RqY4wsL3ksREVx+Lv2KeKuCSp
o9H7bROuMVAoMp6I0/vtVTJWL0edGWAxVISuMuSywiMh2mmALsRrXkac4BfHNXTv1S+XTvlDlbZB
RSbV6Jto8HCr07FzQssCVWzJzP3Z1ZyVEpEgyFrDXBfU1Hcd9fTotauGj8lMoLzR0hQVrsttqzlo
xALLua6cNIPlsiVjY/5lXf9NgVFu8ZieGSfyhfJD7QCMa5Af7tqmNKKK++Lone5MEtJoLu3Z6sPS
Y9zZOIpG6nuWZU1xS9xJ+kFx7b3697dzQ5OcoLRlAE8mLtJWQSsl/4zw/Sq0Am24Q656HAZ5N4qB
Snv4kfF3Fxk7hKgiLFZcHqIoZkAopP9C0It8JFdsJiJd3CTudSC4y7hQEc27K1W+FPUdCDr0BqBy
BRrRMwpi7e4q//ki/17TdCOVNPUbh/aea9KSfoR0MWAJuNE/N+K9k98MLhPB5Egu4lVSruGs7JM9
R9/DbpKvu5HXTHStaLVMjU6o/Oxlo1UAnst9a5MUJ0oRFitr3fTyAK0gUAH4UHmWHXfQhYd7K9ig
8xkWj0Z+YflqWgUUEaUreSn8EASTz7T/l7zxHijHlUye3oote+T1k4p4WkiR2OF7uWmdjbrgTPJX
HbfEAbxzmsIpYiX9iRWbn3kCehmrC02ECRDCY4wVe47/5lxRXCBsbNiZ9ut5trxWDMxlwcJ9EayV
RSykapU0CItCDP6c8oIyu4OcLM3KWD0ggVv5A+aEZtu+MPPNzvwWyU/ACfHDP0vwFEP7tQA6y44b
Dm59+oVVSLr7Vdv7I1giiBxAdpL4jgjgPBvOzVrochL9l6OalyqNiXXULXmwI5Mz0ozLMwhr8k3J
tsQAkcLLohHE+W+tkE1dgvAAfEInjLqTLchQ2WQsWt71bQqRRfVfDtgtqnfpcm0MQUs91NuCZDdG
RU3sQE/HJjr4LFOzCh7/l1jl32ia+fuHQblwq4/Iy+yEUaOmzq995xTFj1Zh5C2067bUSmtACOr3
qn7D00ilwncj1rTN+NmOQLIBb+V9QLPAbuZYE6awpgyYq2CtbUTKjKHgKP55tR4SPVkGfIQtJQZo
LkYdsGVC6byaKAXvI2K0M560RkIrU0J0YVrMdXh/eiM0SX63eUUE1ZBXcII20dCpczFsMo7W7Ob3
TY4pXFXk3n6uss1Fbgph/ASmkOG3xrnswUlhUB9ulpSVE1Icf1uQgzHDsE8COm/8gYVcXZ9DYgVn
1Q4H560DSV+ogRaqDfX9wKEkDTkXpdWl++JHIRR4NqQuayR845eI6bDDHWPStkzbido7Y1Lbg834
WgV3X52kmBQr+7ShiTBrvplosW5xMD24HG7EmCGarnklPGt+ISTNIv5UNXowGcQILswK72tONah5
ERKcZg11aDgfsHQUXjlcDFmZSy9LYAd5aonn03b1cP7IdeiSqRicjDlzf+2md8TjZEFqeqrDQSgg
IZ9tpXW9/gvsDCRIRHfok9OSZnoQoUfiwCUblIixclcxioXal64s55D2vvJvR6QEh1MqN/LIHwt3
Qq+lLhIdZDU4Xzlj94Sy6FdtdZgwMoTxMGeu0VtL7XJY+y9qj2Y/x2XOKhBAJhG3aa2nAH/5Cplk
PziU8rBs8lFsrSlTXBA849q7bdQmM5VFw0h+SBuly7hRv/6fEYQHvZkq0gunicL6iB/sjIO1LZP2
B5SHvAnxAGmR3IT8gAuHF8wbfmd975FFjmDmNo06aFmL7TFYE5wLK+CFkH025iGgoZXt8QEg3uyj
fL/MDHLmkV3166uPdBRg2wzaSolYSn4XbJsmnfpIYTY4J3hX3TjcfLPYGU3WrtXPOQJTpPNMD/TU
P6WFWKgPstinP1/cTNRpfvXsRpapAbARRuhf78PO/85yiA/6TNT5mVqvMPbfS28PR9UhritGWdML
ai2TkW/dhGLmrv5fUblZgVatn8PRkqogEV2DV+4jH3bjxbyeYSCxTCy5pUyJDu4FHLQZ6m0JUjW3
pyodqth+hzAh1avxLj/c0iHIg1XNz40Wh+VuN7usJEooxx8jUBHQfFkiyB8m0TDO1O8HQL5bqssa
lMVlaDAwLialJe6qGBCzfAX8jO+52N3JVzuPkW9+LHhaj7bQ3oGKsvlSjoZaOsfhZKcXlcBFG25f
BGCOuKOkdDoY+ACX+v2oqH64wx1ao8SbA1QzEtcr+pKKL+jyCA4XRYzO3gk93P5Lq2UfFsHu3Lfv
pSz6NrpS3S1/tjiMWqJY+2a5f6xWTNsj6qj9jse7R2auRxI5sW9ljUvAenFss09mbc6I7/kDemDk
ilT6HKdxybTi2s4N6xGxG9QiHJktU3AZ+TxeF6Qfdcz1uJuA/hdU3XZO//XeFCZL/5wwdZnDTYrU
rK+4s/FS9YrOEDHZi6auxyXcR7MZPu+9YbyYrmoQKepL47VG0fA36SviRBeBlPLkLSxyKe1QzmVb
xaKOr8Ior3QHtLsXZIAdVoJMKFloFXRGEy6dHRHiPfagIKaPEiKLqQuuGhh2UvKbyqkn8naPTeYF
FpwTRjBTSow9EEF+xgqHoHLvIofyU9M+Atv1rdIAXDG/OiKpxx2H1ZY0Y1f99k0WtFE/I3Zdp+Uj
BJg1nLjHplcBOqmwYt4Zgh15jdSqhIBxjQBpaanBRo7+ST+tAl8l6Usv86hOIASuBqdfazQgwDmu
BhsuxSlY3bpMv5pRfODkJJ5mXBJp54o4XTxOexzglI2b/+IYdYHpmFExW08Mrq9ZTWQrpq7tNADA
XeiHUH0RWQpgcMTAh3nfBzAjMzWJLAdilPwxce+7w9kRaVtCOs/BLRId63VzetHJ3VoYBYIE/kf1
tiOECaKvzMgtqmdDV9r/dmvMOKFsYAHeJzhkE1zqnor6T1dAmamC70m2MhpIGX4yy5Ttfir5gHXj
8bBK8BGP2KhUBNs3BFAJS1jOWxgHIduDdrPW6gSAEWv+E1AARQ5YKFWVffOhiGBtFYY70BzZVcWd
IGL0DHlndGfQY+4KtbEc6KfSLwXbrRf/ldNY+RIdW/ZEOu2+0P41WGKvZTuS+x7NQdkB0k+FIALg
fRkzin8n4EgS1dp87rP9a6ztlt1sqn5QuHzgBDUAn88a1QwVxtV9ZuvKxPTTsFDX9WyZDyXjCFI7
MYe4G6qpv491uMINwvJp4NvHfODw/135h16p7XVFb+H9y0uAhlR6mRLnHIt3M1dW9Uj5pl0lFErc
3Tf9UOZCyix/GAqhuBrsL6xrS04JVEh2GE+724fct0p9QUhhatGWexcElvvkKzlk4LGG4h6GZcPJ
MHGOD08Tt2UDEWqHv1Cf+FaEInMSbvkr3HE6Q5f0IuYJ0MUjmCsqKnVv1gWzsffZOrgQnAL5d5Oc
VYL6efr7sOuUJUKEGbdgLB1Gs/19ExLVZqtReWnxiDsgzEScCLp5uxTbQgdizKOA+1DI3kmmT4el
UdhHxFCT/gltDUEpIjay++YdMft/Lkky056owRsv3CPhnF2y80HCOYE9DeeImV+9MvL7s7xhvN1/
+1ua5nzfpwVwqFX8N4QwlHWZJtr9TMuV8FT/ZhZsUgd4oO8S5V7N4rb6xAxocym/Os0wUxvAInfG
XcZxh+VfA336gsCk2GjTCP15CGPc0uDB89MKFXbQf2d9e+dBS35fCEjo3pXuO/o8BkQeRvGeb+8g
xiaYz4dxefD8D7rV8NWsy60zfPV+irT0vas7MCFhq6cCcLXtvbGfdUkbnveVRwfbD+MKYmZL0Rei
l7nUMnWlCvAaVjBT1ZFz0y6Vzasitz/JaBs+JHsYPe3Vz2F/FVh9YiTgYJ20ZFPRjOeJxQh0vL8j
faEWPcrPgq5yKWwPAHMGYDYzMQueR9Ytjh6N4Vj1KJFP3Y0160JSJOt1l3QqUWSTkVdYfLXRSkQl
+uPasb5SFOjqhExyhYtOXGFOjRDcfNUzCTJtntEtbMSiMIEn/tLNBf2Lz0In+YMm0JF/oAuIK899
CYWo/PeJAW1XWQH5LqVLG9TLV4DKnCNTga0+Z04FKFgVzTnCTxeh+t84lVXja8ugiwZoi2KjqJan
F5gkhAuzC1R2WiIRP4IOXnZwxQ97Jb87lrwr84slP8Btxd+IxdfmU/P4jC0AthpGIKNUoLDZfVFq
eATSnqwGksv7yG+W6kV50D+u2LwNbmF6qcdODcoQF0C5yB2lJ8cPslRmoWCoJBZvIZGU+QILtmD2
LpeNZrvcl2qaYAw7yqf88sPlKYyEFX5wTuBpz+EffHgnOS2lsuh4CMzKWddrZUndtstM57TUsJVD
/T547rMmX/QKQ3mrByR5s+r3u+mJ5T4fFnFQntdthrTDCgjNnb9I5G/gtUIs8ftCvta9Z5h8Q4Zt
YasHw0x6lTHlTCf+CuHm/hU5PhpFTMLZEU9HZzmCo/aDzpAZeK3/7fzSC6C2AxH+Yw6WXZ1KZtLV
wQNYeOL3BrFO2M9Tc2FtaZvESIyGqJxKarn/YBt9etbdlAftrl+zGnfq+ffOHhFq50q6UQJEeB6G
mKA91rwFH5etvXdrl/ZCSH2VxXD0LPpGmFu9BaT6fdiZx8oqHsr38uV4JsPhWhCYLmn2LJIRmIYw
no8PLjcW4G0oAPAewPOh3ct2QQPZsoQvQaEYBxe/srdrMFo77opmjqm7qAMe9DFg+US9iM0bjDiS
ujMsN3IkUho89RSGZwJmPo/ZWnF+wOeGhgC7XOzSRVu2qCuEQe/Y37VyyHt6GwkeJ0NrHJGpotsK
56eGjjnWutlrIyYu/bst9yA87ClC4M7uMpyzgfh0D/DjV3+OspZx7T3mKKU5efhEcimwi40ogSJP
GA/XI6g3LzbH7dsQvGZItYHAu8C1Ws2+1ooM5H+w/HlQHX4mQdyYC1BI2WL3oIheI6r5s7VQXwAo
5YBQ55Ysbk/WmScnZ+aR7SQqQSeJOJnDHWMRxSyqaR+vJYTQQFXzHWQvQ1eyUXXpgklV2VIUuySg
9Szb+0oZWXMoDTiWhEvUaEMSzh2oudfwN6hlNk0BxycpSfwaL7vtVLUEUFAFX/hTJzKwL9a4v6DQ
ohthTPTFyO7O2VuKTNiwoDcc7usVVJtNIBclzGKighhz2rs3toLYM/HU6s8TH5aG2E8/v+np1EQX
5EUqIKWBVv8DF+ekEUK/oNI0+9NGy0THy5xqinlhCE/806W9TDhN5Vo9cHVc7sUTvWNyp+RvjM1R
prcZt4eAb8RjiOTeh5TZljJ02xKXZ8NaRwjId6usg+4niPtm9fM7ytEL9jQEsIE1Dp3t2F3cgT/c
bqRFtCHOr4Vlj0YucqZfmSMzdy6PbNz2AkGNy+C3KxNZLTYSX5k5GgBc/m4qbsa9rWFLNARrcwaW
dCkL3tQFQWAzN4/QNtUsTEmVab5p/tR1YZZsKCNEZ0aAnZZZHW9j0WORqmyh0psIEou9CDAnDzeF
1JYee6LGSr++yG2NZ4DbEe6lDHH06Dwpj24ZUq5x7nlXMlclZv57HhU1ueZfB0+QTN6WjpO7cUnu
XWSN0Tmzo/Io+QpdSr66HCKiLEuSiPMQeGPVwBE86HLLce6ePtQMYI4e6Jq+QZQ3HeJRgYLSqVXu
qDEcRDUCSA5mBfGhTpbQ6ojirWGPaMhhS116uC28L0iuxfofnN5gIPeM/ETMdTHeqF7B6V2tQGd8
9scPnBFWUeOec9e5iHpIjkxccenu4vfPp7Ypo7NlsKKVfsPxSEjfPxyXnLn3/X8ruRKwn527SsXm
QHAK14mzFUHHn7G8OCtl4gAOw5ycKyrkT1D7+shD5SOybT7RbD7y+GOIGiuSsOwNNCXUihP7Uu94
furjOIdAkn63mkv/YrfQu3kg45hfY95QpTkpbTLI+ughU5MKAyc0ZMGQF65ohC/GHd0VaZfB7juW
iZHWBqJuLg+qz/uLGC1D41s3EIc6XnKObe23P1jA9QgRUsU7xgskdxZBXHY561o2PrJERsUTUOyI
pFVpHiNy49hT5ARH2cs9r8ccO1FBzsU7MR84iua0aV+RB84vWaIwMVlm3Rb0NHoPOcK9J51fmLF3
EUdP7oKg7KcJmxVVq2Pug1SuWVUela0pp7D86JrCtd3gG4CqmNWcdMTqDi00VekVcmNDNrre7AGK
fyyTDdOsbjBh6jtF9fTPS7sM05Pjlus1izD3r4J/AZ3pCnIV/en9pL9qwxDOSuejlghJyVcsmzW2
VLuHz69j6cpq+8Go7wDpB2/oeJwDCj0Oiln//klezUZghvV8W4001c6d7SdusDaE5NUCMVMZNWl9
a7kVHdG1VHOdsE9jjwh8cmORqKFdllWup8P5M3EVFkBlslyYatJxDKW9MUTimMbL/Cy+Zn+5R7Vj
kLOt9tLEnunL8Q2dNZaFUgKknJFKc1H/iMEyPm9ssp4HZxg+egtty1JP1yFIqmGnSVkUoA+aajg/
/v+ydjbeR5VigDYw81ymHQ4d2sPpU3lwZFNKyKD4dMwXIDOlr4OlNRe/xkIK+VJHEApSVdR5r6B+
j5ExnFuoSGRfjl8C7ySRwJFVXS7c0dH6yVN8pk6ZF51xNrwxf/eTvNW6Pi0l0/vqaH/KR/0omWNv
4hVzYCW0u1qr5OEbdOeJqPaqZ+5lXyaoZwg5tFwKNA/xEZUpZbvOdKZltCqmghyzzBwMhZlvX0r+
sAm1Ek2xhO7q5UI4RnfDAgvjug3/LxJQak6VVHUKcXWODmsKP0oMCTbj59vshg48SgS8A9XxhCaZ
jW+gPRAk+vEVGjPi9gvPRys3ZI/VfsL4utA6VPiWL4Vy1TSy+xRbl/htkF2SxAKW2ga8t2sw/bXy
fo3hTIiMgkYBWqBWAEMObw3U1iHhduiEe0ZPeuBeUXzWk4EeogxAdKi0C+8O+Cp09qTxlVE5iihR
Tdut0OyTaTjUrGwSFLLmibRCZegAfi+4iQWHAqniZvd2ug/VRL10c6s+gjKOSk/DV2b9qveFlTWC
626uAqqiSZmh41+CqI1D/GS56qGQRSQP1qD+oo+dmKWjurKWB5DS627Tbn1lXS3WVXhX3vk77CUv
aOT2WW2/q+aAALJUOtlGOKOS9TehCXiRXf9JLadHQAf1xWCwb1P2w2My8+xb+8ArzeiBiQ3W8Hd/
4DJsVT6IEquQYK1DXd9ldsB7OXuTfWTkQAIL7y1umLHU/vuzIJWMPXoOeg3PW1Qm1DA09rk42+Qj
n2WsekS9WbLzrc6rT8YZtUbl9G5WMOZf+/7G4TZl9DKubAnWWECmMJkQWwSK5vOyatOIyDT0ET78
Hwh0Xq/XVWsyhxfn3GdqLdp6NNN3lXK1a8nd0DwFwkbp13L6o82aKiZ5g+BMVJ7+iRnrUcacy/G5
XAlkBorqDGXBJyK4w0QyicKAMXVh352581PcvBfTv38+uVA/VTOg7Hd1mzj1iJus/IUxdHtBhcQr
UTUZpmzMApbDbr36Iwy84RwfoFNOzAX5cwInJOkSvHh5y90108Ppy1CfF2bOlCcFthb6lo74g5BM
uqKab1fUMoOn5L1TM/GqUpuid31POXY+ItmTj7O8LKAZ+3FUTxCx/Op1m5w+gEqowD9XqTXqpTZp
9RoItDicpjv1SkDaWAisboALxNG2jt3p+6mgscHTHH4k7mRtyeC1mUM8gb4VKK64bbQAHuryNwOh
hsgV8AgZ/lrVEyQDQ3q/mJJLmXvjQxIMfgi3GR2ZJ5LDwpyPXmJcfJF5h0rlMLFQPjabBNYKYvGA
P5GoMN0dHONgH+8A/nvyPyao7lFWPlOJ2vPN2M9QaXhuKgL6RpzMQdLIvwva2vnRI+2Jdg5CmNPp
LBJnCLPTkIY+rUl8MHVQaZuPch2G/Z9oqCU2u1hyhL0Vc3ZS+v4tMLpzdg/KmL5FJt0j/fYzaa5v
QkU34DjugtKnhRk1zQZ3QWEYe0asEpkDI2RELfz4nRUM19XwgQ0V8v0znzmeWNHnecgefWQ+EJQY
IPFGGOlGLgcUhdDlm6Amnmh7sY2m7fUC/F6cZoAUk+1Mp+F0ucCKIDJi7hsSB05BVyzVjZzrD7bY
JUFcqjo2iHBWcwZzuPX3nfn9rGajE90H1pCDCn6d0A9v3myAquBH/MdZDUQtmSYchlAXDPi1Fnla
t9jYivJ7WGroRrjx9NI5U2E+OFRbEueNWhlOf0nJbC+ZOSf+xSinb1zNl3kbHmyoz9OeaOA6+J30
RiWBFHAJ/li1nABwkK+AXaTxzJky0m3ejCl01AQ+93GnO1yUlOLVPOZwoctcFpJTGY14OrNkb03Y
30wyFYOayiKga/cnNhr7OSbo3cXXGPp4PHnB5qlada4Rvqo5z2ZleM03xZOnU76fakFpnxrySag9
KBGb8uaINDLI6lrnR58YiJKYem5lkFB50yJmFi+1o9kbS86Xoy1C0t0H3ieZNJOww+sG7G9tG9tG
2uszX/cf06EQaxjRNJuvMMM+G5WfSGDWRVdkrUpznU3vCIWMthZjE7YM7nMZ1BKszT2IbD3T2DZF
56SANPnS0kWTATYWs1E0vQAZ3Nh+CTVz42JTa89gDdVZWBjqlcPqyJdCAOR+McuM632QeGleGExo
njIPAbmqHdiEyOmD7AcVHA6pnZffJg9tSwiot2ak4Ih+pZirKOM3iL0iWgxpy/RUF9t1fFM8Tfzk
f7xgdv9LULL1ik2PHCqypU9RBkfIrtTN2WsXjJDtoFlmYXDTDzJLSXgPeXbaXAyuSEmX7jkkqA7E
h1gEKz/OVCNa+MC90Ds+94fCVVdvZikncf2yF+PncM8uUb1LlbeeffJuK+FWrahe6l61LVzEm9My
yc0zjgLsb1rGdsqW3ownm9mG7cQDp5b0ho7fgtP6M8emwR1ws/ZaljoE8A1XUqUQ+x3cyIV45NPq
UNYVIKHfNeEBBoIAUzaN/3mJIDLNrhXGEg2EFoylsToOS+u/NRyIYB6QltcEHhlXGlQC30r0vl9B
vRPkqKNscL29FhiPB6PAnQEJPQcIrX9+0lQvYbxFxVTjdcpEV0yqGyNSBIUqD54i2JF9ddFATWAC
q8EZyIz/uyL0OU6LviGW75u3xboU6J27Rp+svX9aNjS9JQyG4ha1RhpPwnyilAYD8ZUFdz2l8pWE
Efhbki6jHmfCR4GsVLOLA+869Ec8LXUP/unUJQPg6Q/OB97waYYL1tpPUCUxOefhBrbh+8p+tUi6
+4hxaXD+OwY/U8fcU1CEhwMZSPFyQZuT2fNimBp+Bo3xkOEN6sfQ+Ux33X7P2McGZTTpnTAyQC4w
sBYxeS7aYpvi4MGnkKvDASvdWItAk/zTu4UTkogTrCLhguoEG6lUKxiJs9RPGIYPB5O20Lnq5r3+
WhvfiY0E3VzB9nU0vZv/Q6Uy9Pot6vZ2Mr1mFCpqbZbZjH18t/g3vayNiu11SKUfMMccOW4xvPT+
CkQCJ5DRWPDs9uRcvfyDKesJWMp0dI//S2KZwlbWHE3ojE1RU0so4Tc84BfSb/dL0opYBxhRYGAg
v0/rz9lLXSkzZb0RWpV+UMg8t4UydB6CEuWgRBnzJHHC1dGPqfB9BwTr3a5CFPHPdlP8SlpFIEnC
nz+e19LgNHd/rn8mFG+zt3Vq/tw9fvStxqNyvcv71M5yXgcNV2fcIGBbA9xufWm+cnseVOOCIfuQ
AyQNbyWxeTat92ItXaTqAcvTOyiGnZoN/D8k5C/eMv9bxLAE9l11qiowyb1yoIFTb4MpaFgcTP36
vy/NydoxaFYM4hmBYM0uWhfR88bpJRnjqgzL7uXvLr9nd68F1HSoZAPBbyyyQrNDOcxWqgG8yOh+
U2bddLNBlN9xy9PERuJRuHXNtTbCUS/yOdO/EkBPJlFtWK3Zy+5hy9DitF3jnJhfcse4OzJToPHJ
ri9SPALZ546p5M+LpIgsswPEnV2N+Wm35+k7+j5zQLcGy4aSLhyD3UFtCXIm3GYJsHrR1biD2+qi
ou2Lstjl34EBSIhsqjarZQ5v1sMgk2CkJ/4CH1CbW0KN+0/UswN21y0ZdmZ7iK0F/aPuj/wGgDLf
IiUvB5v1aR3V3t/id2qGw7maH5hYLxQe2JIPXHoPHOSn/pb01vYqbQKmLGczUBxANh+8vkxfpQZR
2DGp7/kr3s+qba5FVS5dDhaexiaE6SMoa4n5IOCcM49qTdlwmtBVLFYuprbyw3ivjDq/m/FU6Jh/
u/ipZTTtmWjsQ4szKKyGVAGY9ubSxO5EOIOAqeHvVs5poNbYbGOm+0AxaxFvALr7DYLzWBJpWEY3
F8aMeOE/cvkXZtTqaHZVr66IXgODdXUWTyBK+BBD9jxMwjvLToCuaj41CGNtWex3fWnNZLb+nIqK
7sYqcl+MxWGPpuC0II/pg2teU2oOqjw5dTj3dtMjs7RAZM/pvNP9MXXOzvlOInpvcYSw4HUWemgA
nLNLBFntm4OT69J/hmCrlz3ge0iL5aXf4aq/g+4F4WIoxfZ+Qz13DDEUjnENFwiqwS+3VHRrNwRf
DU1zfng2dM9UOTZzhKBGVl6Nz2fWevmAjTXIBTYepe6T8ZtJaTZZfEUZArfF6qV/UgBMf029SeVc
SIJYPR1kyIoFS3/rD9IQwyIApwWng0RuPo5U4R2C7W+3jrue1vIPCRYBIJtc2zHY4TSV3sVSUOq7
oU9A2XQQ/8FkFATmcG1vr19FOQXfGhnS7bUfNqG0jAk/gCBfxMfUehAHHVhZTmUWxXNrCNmR0o4+
7vu7sWzkKcSXNd66TmubqMU6jp6DDCBxHB+fcIbZttHPN2d6PaCUKWN8zqpVpQE40zszslrBbYA1
sjg/0C5jWdJVmYmvHWVbDKMJGf5aR620KITTom3ObsrFAAKzkEGvXI1HOCyiB6bZreXaUCmPwNHU
ljUxtCqxy3UX5s8CDtFa1goGbqgGuL+XV8rjwjLZ4bpcEo/fcy5yYTgVq6HvFypq53o+Y7pEq0mW
sVwHFpV1vQnMg/wTvMukvs0XmAoEJ99WhMMKdO6JhPOaOopKax+keLGQ3brf5HfGL2uB5XttFVOU
KR+88nKcX70yj1Gp7FLxJH8J6hHJZk8DyOZTAmPeoAVOa+LK0HuMqjBWcQ8e0zf/vaFvfSvmi5zo
AGgbz0sRfjWOZV9n+HxCx+c4+daBnIKg+plpPdLfNb5hLDlN3ktyZW/as+cWu2SMstJLlKzkrycf
stvZeiiZVif4SZh8HAq1d4seGnq2pb0dr4E9Ic/bV0UVR9qF4HamDp0DCszc7iKgkI55PbaxVqP8
ccY+fk+Pf9ZjOwvrIRzwY/dnMEnuUKFkM4TkVIC8LXxWCpVAcQ0vkxMf8Qai7xETdYMGR/x6fH1C
sgkQnUHj9YyHppAhB2VxOAAxAtjNl/h+XQo7qwtL3u2lizvWnpolEIeKdtdiPXVwb5I+/pmSPAkq
a11S04eqMNxX2GmRuZ0dNygb8ZJNcq079cmSuB3+Galk8Xqp2lJmwKji88F6rKL5jKGKpsMUAGuU
HjnMyxcxlmY07ANRsBUPF4LUa9fYHpHGC3mJTjBBtSOzhzVRNPsK6gKVe+aa5vincKp7ZsOz/laO
HSCbLnpSsuuSs8Pe0H/sSH8CiDAurl0X/HotaxOBYPzZZQQv/t8D31RCyBHFqE3LYAbmU9hNmk7o
lECe/o/Ki0aPB+LAu7cq7bQ+9lxuRt9Hg7NeJuTg3i592vEXg+3pbcN+lTvq3jQg1Xl9uSlU+brz
dcXrzzB3cHZuvp5DfmxM4g6+JbK2t1Teeqbe+sW2r9qP4BYYtNB+RF7dz/9na+YIRSsC6WUDsGeL
HPo6NDLFsjhBxmR1gpveolj53x8aNpLBFHzoxzb1ifmv/RZiPVLVwTXvr6H3EkEpmC1wX2JV9UFQ
M2LbfsUTXpuVEYujBkOvknxBiXNWTnJbh45pjkFTUhM/GpUqt1gNZPwpPC4KRMStZ12lckPavA6O
fDImWaq/w3OlbaJCMhUNuhqgy37KF2VhsRqZI5x8bEssL4GLn+qtPkN2PbqD91RPV1vzvnkKSDyC
4IRemhykawk5vCBXvNBGpB9YpzgTiBEUBxxb8y9RGXWOVb/07VLfNUgkCseuQ+Vf5KjyL6TVptQy
A4LmwhNbaJjrL6NKK4gAq79wweMhC5pSUluG3o9atYzHJS+RRp3EFCjtmM68kUi1MFC7F4B27pWC
yZptlVPQ+u7mwSqARRe8rerqCUkmGAU0C6wLptNMoUsW7h7lkl66LjQPCEc7b1M0jDhlMUvqXTfh
sWqIPbh7FCDsR798BxlR7RPiPjc6JxQyZVtm+G0vhXmojCAnlPLwbUKriCNFxAX/T6tBx9P4LyTV
IFkpzH5qEjtUfY1Y+FEaKdkhw1DPi2xPCAEtVPpOXUpQg9e1/p7z8kEh3nJySk7Meu7pP+hgJJE6
E0FhxBmM4IV3E8nhOB3pjZ0br6arGaPyppvACR6w4GDYIfzgm3uWqGU+sIl/aQhjdS9V93K1B91v
FDKcTC1ukgf5Tqap0Qr+Z8RMNk8Lg+fOUuebtKRQmPqzr2udbIsLR/6K1h2/K3vCopbR6QRish3V
ohT1dVaFyMyJergqhkU87T7lEIm7fyHZhOF1oyw7oTzQE2g4eFq/Ar+Ne/2leSP/v41xk9VjXb1q
VGl/PBmj5PDBE2et96P6aFfSDPTgtxlWx58wYr4pqspLlKYF0gK7dCPh6NNEnn/I9SJ7kxH6MZ6b
o0U6GrSXR/zTl0RiAzaJI5RgDgovgs1UZtfwQM2CYsh5e3EZaOizq10HmWfD8nL2RuZkYBzUjlcK
1ZT9zjOpo1scgYzHdfT/icvON003YqtkHdB0PjABDPW9WRYNE+tX6foNkV1LfYibbvqCCHtJoCMk
CUkKNeR6M2iAFACm5Oi+SNvaLnfyQ1WCcM/GOCnQ/jcwsZ8cN0ceyt/XMqsfM3AvCYKIRUKpH59y
9Utae/s0aHDUXCdjPwcKwDXuJI6G/KfmyK+E0DZu7aIFDI5CZI8JVWy8/QNG4Zgv95dqIrx7x413
LiOdQbJj5WOVyJLcHUDMxRrhdD/8cjR4YaRS76gOmVxxzUO/Kcq8CqMb7r9S528IkOOkoHLdb8Ux
8uAJxoqGXCQCTBFsLRecQKRXryojnoOQ2wS2nivuWKMKXYY8CTCXZlTWwKrbz6o7AsylONKUaqv/
dTa0K9EoehBglKeBG82slL7qoHbWE9LtiJ+MQ7QGzZPvMWRzoS7M/FlOP5F6kHMO6Q2bXfgb286q
Ae+Cxy02SvQXqVlny6gD004R5JUyqXkKyYJSXS1x5ltxOD5Oi40EzasX3ByKn6zwu2vbx/lxlHEG
cM8nogo9ez41oPw2lYvT3Cb2DJpkojvIOq9RzGi9clqYi07Ig1xtDLTAep6rRAEsBUjYgil5xPNS
az8gIHXhWt2/PRZTYzq4KI99Y5TO8CexamyLkGk9HcE5UNqlndxY6OMSaMCfW3ea6yx3yi2p3zVv
yzkIQhBrGLdG9M8EGqXWoq9RTUuesRIWqo47fMM7C3PV/4m8s6yeJuCL40FzvAicRxIK4CKNm98u
nG2jKoQ4ZEtcW0TZqPBT4rYMNtLKmfZUIGh6bMARbSq4ntnEMtBIK3+wrW29JVp9bMDVYWlwZqCG
roFmAIEgFZwzNbIoGSz2FCrXocj7aao6kOSZ89MhqMSANhgHP2dXZphLDhpUbtTrOJKHaBo8Ymyx
EYrGEoS3t0WAu1MKjajFxfFAs4AdmupD8LNaGZ+Dfyv1f1/R0s8MwPxjLVCrRqnjgeQOXei4ETcO
nLMtUQofPepcTuZmpzQFnshKkE2/hT88fzY2FrtTKwyn/IrJxSpwa3OTOo58P08hdCwzJ8mj1E4c
FFYGskd0dDxJg1VZbV0LdI+K3AZSnsiIOZz6rK9diMPeWdUdgm+ZLHa1WW4DOzwwC39DQ4BZQI8j
0Ryi65A250OvzR4U4LVEMPNqgVwwnwlppIxiypjL1cG6e0jCrYnUBfmfcTt6xUBsQ6Zf321gv3tz
4SV33YVHrxbRoogI8feqRrlSCETLJaCh38YX3m2wXD9V8qpS+1LS+AOvPF09nHc5JXuPlDRM2SrP
gcdjx027joGr0jYHZ4+0+FBrDlK5xCvnhbJXEOGFk5dpSY+CTtaso8nu17YOp6JbvcNVsHtqDsC2
yJVOExqulquI/51n1eWebA3ENQW3F4U30wARNw4xhZe4Ax9XVo2BZlJG2Uu3sUT1mhBHkz4n7IX4
piDHVqi/fdbD1cIEpS1FG0CeAXK0WEHPnv4/6g1KnQtRGlDwZnUqFlN4t7KzGE+99+QbbslopZ9l
0tQwK1p17OOwpVGfGudK7Q3FaPQtbuUmjrQdsZJ21sLxFyr22THjxRvG2sPI0H5KJX4lE9eH+XAM
XxQ94aGDHGpGr8D/TrO8jlaQYeRsuWsDfpKQ6Uk8iQjlXjj4tID0jhpXg+M3dyAJrGU8Hg7eect/
Mmei0Z/1hNbc/QV7FYOyK4z9LDOhJgp9hy3elfumtc7meN+6jffM7qpZ81Kk6ANWS0StLtlovNmH
Se4suiioIgl3PCs+FpHs1EB3w9VqhjVaSIVRZdMPuelJcxWpt7AIaHxvwKQfT7JAeyC+dnZ/G1MW
kPYkj7N80Zhl/dsVYlxYNDr3dCg1PlppF1RyXI1792jiTlmDaCMVWnro2EvoA7g5REB+IBU01xQY
dIGL8jpDnA76y/QuFsKGcddnIwyURQgenTmP4DXb1JERhCrXw4QpYOVSy4HUPclB+4xxpHIpgPCi
8yO37Db9MRztqsOnjTY4M7ZPeZCInHuM0+EYuwjtRlYytVDKFPXDuTMacos4uPXLpZObmVKfrglS
YkTi8+aTHhKfEf6XJmzAsmHrcO09eHSu0EDbCw7PorDYrvbLKhwIRWHcQHNNCtdyOrKPca+C4vp/
1+2mihtKvrC8245E5jh89ImfJJOHCOXZ9jibCCE5tIGG5RdBZ1jidsDJUPUh3lUi9+HyexAWjFFt
4zHSFpBTR6KPC2MwJkJ6NgUMTAihZv/lb/WBkQ6n0N4xt3mHNAhsh9fFwr0HRK65g+zXBnTSULQF
G2rzK9k8zyfHtYgxC1jLEJHI4QxYimxzq/yc0AeoQvdxHzK60nHjOCiX3z8PGIVllzVuKpPlhVNI
drBkxCE2oE4VSqFKp+2eUttCJs7HnCTrtbk4VWmGOTORroGTt7iB2bZtfd/VBlLgf+JlZiJkLocY
W9bwFU5oaSbKarxo7ch18ljejryJB5rg8CHDxwhv4iuiNYWYcTynKPk3yALSP8WpDeJeWHHKpVRQ
VGaPcbNezsTCTeghAPVm7JbGriXmeyW5lB0ahWipkVAfNzLoE0IN9+J6EoBgRaRwXRfQ9tCBF7HA
cgJZK5uw97+uqnYKJ0xEK9BpICafErJyJdEQNw7JGfXgbPSb6yaMZ4XGyR4Y4f6MU4AJxO0q4O15
vuDkYYWdTKlPgiOqmmr4SuUNfvqLLNgb8nF56XpbuNWzL/PIMBL+XgKjAV31ShZRqwUXaOuNiYED
5Qkjs7poK9vAtdMQdSHWwxpic+h/ZQmLiOZWcK6uWbPK2IoU0534tuu/NGe2NM3TzGQPT1hl64V7
SMiMvJgw3WogbEhV53n6nrDvg8hgo0tR62fEcM2+a5iNmED9omPrPOBnAHm9LZnrLfXf7C/qwuAN
MM8fKHiWgMpFPvNcbu0iV2zppfuzm8O+6WB5INyFD5Xl2itLj/sWlyPWDQGqzpuUmxEqtya9LK+7
7DWlVttayu75/l6QmLyGzafcYlid7/fvVBhj4MP9UkGJTn2Xky1yRh2C9jVrLUAHaiCAWhR8VDLM
hoASG66aHzk2Bzoy/mEXCheyotP2uazlr9GiGnj9uHQXaef7VDJqqUukVoPZYQep0CROJnpQT8F+
r3fnaSH7zJHEdfGibcg9Sbhdrs1PyvKkgrvRbCS+gxp/IurbW9P+naB/k3z6RdahQoCp3GiZPfEf
dxgDf4ICnzwtPkiPSfpeV6UAlQWXhoYWhwvKZ5jinDqpX9PUtYIehAuS+sIVhxdpbthYPIVlv3o4
sWe4gyN8AS7DMmhCZdlE50wnVeRR3qoOIcdOvVoOGMGPF/yY/t8QtMgbhcpsecAz+fkKPZKbpLON
3PQzOPnf/uA0uFSXLT7S09E5hIEjjFpTWn3NcGiBC+1Dz+ipa0B+ngtdJwD7v0mIH5AGDn5i65S7
5vkp8BikK52Wbyswazld1HlKa48kAfqjrc9S1MzOsO57lr5J2/jtlKpMnmdy5lUcNppPJET/jtco
xbxwnVz7Y6EY34FWfxX8tMmW3VfuiSBgLSvORancAntEaW1d4pRXskwirqnlVHfqvo9AMv/EWdF5
vp4doSbUz5RVnfLtp2wnD3sHIWxc8Y7Ka2tppz6/4eUZCX1kWVAglS2QH20+BBJWQLsnWwfyIn0g
bbqiOtt73CyA9imMQw3AZTiWURgNvcop6txT62TeMYG/+h7bTf0pjMH/IfcKw7cjafZyhNTKZydx
9lSeKDtdmugfMLtM7z/n+7NwTtrf/8NbgdpcbeIBljZZH7Dcoz/5bKUYmbv78FjfO066avCvwjDq
VqGuVxG2j3TtCmaY2PnhaOkZy4ILuBRtAS0oW70YFqNT/vjTEP4PkkYvBwr5Xd6L80HPW1EAuUjk
XJfc4nIWQWl5c9PnzByVs0LSLEuDHK10H3ceRM/Qdo5lAwLm8SWtzDr+d9VNtWTJbPMrykChFxPi
KV4/cSEgg1tbARpmC/fvvKAPY3sxI2Qvc9H7kKL36z26pqOsAZstxP26MhbDOdqx1PrscrxiWWAk
qACKVzcXNhWmiD3zpICRSg6tfoDyt5dxSOcd9618q5dM8mKA5/R5ZVIaFJcIU4rmPbY6nRpbpeVr
OBlpwJL3gwRqXYcdzLtGAvSHdarWTyNSVH4DT8uMy0byS1kGQC/8CkrLc3CzhGKzzZkxZgR4UVdx
eY2aW+wjYPy2+xL1FS4RnV8eHE90INUj6505U2hfSywBD3JR7l+LAannNIA/a/zWVBMQwfzTocIG
2EEE+Zy7IGL2R0UyA723LicUtdpkgWj6FfGEpXKhIKPps5BiHIwFPA7DuNiVzleIC0EAYVpmBABC
oTysIXaORPYxB/uJcwjRsF+AMxl/xflEmK4l/UGtRf6/tuxqkl9jfIcrskADp0YGGjY9DwiFflru
QRWxw87rfYpN7/0kEtNLKNAv7oEKEyrIPg1a7rjnKdVkpxBSkCfK3QseBK8MW/e6o/aaJ8S+IQuK
VvW25NNcZ+ubqnuQiXaE0YaNSh3bdKi4Q5xGrtn8JQIcOqNrORykYP0WVpKg5DoEbOLACiJOqU7Y
Y4q4EHYTdpf8WU8TqzUx5v2DkJmjrkeJTqFOaELYOmzYYx8gen8rHEvdkO95O6Fx+IRSVsoDDo08
L8xd9j30OPxIknapNJOGCRDTB64yuNxHx2P0pdFyMuWlrfdwqQntvlawjeb3DtuBsymlNFnSopa+
z4KdEs2v/OLocfVXM1EINpvvmbz3AOZUGWoybRfwK13VHHDo3JYTQsg8fvwrS6kCQW7CZh6Tpqpz
QlTzyo4dGU2bQdNQlptpPH49JeCcUhXA9iR+tfaoul+7i9pgLTk9k5zmrRPmowSmhuNfc9CU9WtI
sM6UY+yw82AF8E7ru/+dAFAX7MELkcrAIZkHhuF8T5q5Q2lEmtg0Smym70wChMH/B59ih+0lS3z5
7AMz57YU057TFGBD5RW2QI45Dwz84JuN7hTDDttYwUWvp3Wwkk/ZedN3XDKKvi0WTFUOdc0Q56ym
6qFP5wI/u4fByA0HFBnAIMbuBfXp0TyhheauVxQ624NZWBAR9gop17yRcSzHRLQieSS3GF+PHAj6
bE9cwZ/onQ0TcLMrahJHGgL+6F16/37AC4/TEadh6d8AksOh/KrCUfF5ImRBiaHErnn2+lhw/8hi
h2AQIUB5cVgKy305UXkw7Bj4e3+gccdj1XGGRvtXSRWZhyaLDIAFFgOgZzbJOOCd55xlSGS10vJ3
5uaTyVDj8EbYHV+BtjhLEbPQd2SI2qfeETvkrTzIz2V6+kZjUUgBpOjpDtXbaMplKkPUL/bSMYHp
GHeEr+a7pvutCYSiek/KKN4rmAgCA8f91FId71Aaf1nLEiggtxIFEC3CMvfK1zx3DImmt+4bVpug
5fcp/cv2kCBw2rszVXpbKdy6nUWUI2M+nRm7WOpb5xHwUuJBEJQqud+iLlynPsw6pQFfi3ZV37Ki
l5r2RIIiVyJ9oRZauaYfWoYqrF4RkZ8sydtahN8TYXd7ql7bpUrVyNNc/moCdfUcPapw0sCoQHrM
WUGruJSn1f5PEj1++CQ2J7AnDvayNLVB3O9LjoU/o+ORZS25i3BgO2+S+n/iZK08zBgcRF1zoWdi
cOu16/HnuDEmsEdlouS3jRty34XApO02JEEPKe7vKxe4fCCR5etL5LhPA02u/FcVwlhTu090+neD
BVPmX0+dVi1fEbTAAtMKWPrErocjMzrUutD8vMyM/qBH/grIZAIXF/mUz4fUX/zRZQJ4He1/92i7
TrCdPCk8FJlU7BWUsOX6KClhDqDfd9ZTSPWSGAeR6DA/nwb5LUcQJQWZh+mpMC7Xfo/9lF3cPtyP
JqGSzH+1wJfkZ7rweUXk5H/zafiNPbh3xCsc9kTKSAC72T8JmovpxKqg9cZXaWwSl9L2HEaiitsi
hPRK9h5Ivs8F/sZT4kNO/4vaqumHpbNvdrVLW/KVjVq/+xDwJPydj7fsYpVsMNyV7yyy+rXeJ2zi
YfNczV2+/Z6Rnrqr5pP/1l9EPGu6kLOh72DXgIb+fB/2FfYIEcLw9bWf5CbSYrYaouuPHK/iF8UO
4oeu9RhuJN9j3xSi//aUaeB70PjdrCLUH4/VFaZbI3zb/gl3rTKwecCLq16PRM51rC7fGn4OUiqz
iPmGy50sg5egOc4c3wcW86fFfmCMMxkzaszrfwKt53BbvfdC4lZasgiBNuBEv6qigqUEfG6K3W21
ooi7Sw4t8WK2L+zMWBStcYE8rBi3D+G9YSj5isAOd1EdZrIKzZC19r3DpattMlbh4768SXQ4D/Ax
MdjM5oiE74lK8Zyba4wD67smz5RbsY5uotoK56e9HH+wOdBbl9KSgToHlx8v9m4NpteQjTsqjYLV
Y80RDeLM7mVhWMcPKwVfEB8oJxaRNkQmxU35qhxFPQ+V5T+ORCjNdSaRSNeS/4+vqU3Pt8uTxUbg
UjtLD2ngAlmhOkAJT2bv1j4UcIXM1n1+ZCNKLYMiQAfJ044SYpuH6xwSLUmryIkvoV4puluGC3Pz
kW5Ekx5DIh6cCi8t416iWJofnQXVrTDZJJBK81+pxSlPRGjaO45tDnr3NEIF8WpNl5z7h5jbtf2p
HRcQAxzYAzDF0aDdar0BWOGdq9beayNvb+pxvLZGXBkqvFz5g+zeNL3tawDvS24dCG6QPg70M/L2
rBj0t0bf1AFPevWaFnr0SlqdqTGWST30S8MDGYf8xrH5A1vaKz1bj8IdRJj/pptQib4pOSjbieEY
piPSOQmXukw1emz6251NNmSGJYY1ECNtvF7zxnKkaw9043Tih7ymPAC837dJOPK3l56sKhK1a5Au
bTm3ycU3n1s8ULYzOJ1C9lMni69Wph8QOpVdyIKpiKkj4RfC9YlAXRE3wueaLWimRkIYQp4Dl3tA
37fk+f8xRQUi3DiCHD4rxoclZ6OICzjvn/ohKFgPBjSuTisipNhMitRjxSXYgtJAqBNsMH3iuOTe
6XFv4gOvxwRUhmQmOgkl5AyGUm+8pKAZHeirQZ/LbgR1GHq1VG7JueSkfKXfwM8D/w/f3fy/mbvo
+RrFQMquRbNuaHgxzJG4lnhOxWB/gdlYTPGVmnEeCl2IRaL/Og070E9KB6OpDVTo+L3XhoaUKm+e
lTua/lunehiGfWMjyLGmLnnEuL5WA5kfQOQHO3IHK9LSM0bj+WIVS3d92GT5Dcm/+V6WPEZIuJQE
MofBsVtMQHfKhV6QKfjSLRSoPItsjtztw93Ij7cKfLp8iHcHFZohTDIggJADG1MjrFd6BkN/1EaA
9L42cRMePT4sB497Qd5aOUMPil9vTVGZnECA3NzveFbiwvmjhjtewJbmdXDzuBtS2IQVNDcSzd7f
zzG8PAkFn/F9awMtPiQ9dfuYKb09b4v1UMlBP0+vdj63R0NavEDc4CCv9mRqSllNIzfQud+6sqH+
tZLk51/Au8AIMlU5ykaM2ysSDSwQ7p9JQ2cEsf2X+EIcuqcTan/nSz6naR38bBnMwYhZbMDSfnPE
DtcUuK9jwxmqD2sihgqKmtv2PFhmBRXW0E0RcPc8Jx9C2A9WY+0OfwbsyeLUx1yUuAs+I/qxVgs5
NNtQrMa36G/wGU6lKKoTrYhKdHdcKVv2iPPmpBLfFZ6km8+Pa82Vx2meaYsZGeEhzywlPYZANFjV
HdKq1EF1U52naf6D9X6tiIYGBAG5J0Foc/0poLKLyLnN7bQXYR7DD6PDsqmI68I3cxO5A0QtghVL
3K0tjK63g6vG6uZYTMN3HPpifX0gphLEuVu4Vwi6y8WssUxCBS51czC2PMPPa+BsdGOJe7+GQ1QK
DVLdIONFs//SDQbQwsROVqm1TBYqwITHxJGf0oTOuv7bZwOI91lvY39LQ+y1PZNtS7THDJNGkA0i
E8II5U9F9s1GC7S8u8ZrMqdwrfSNctAIwjDdBSyutfIg48Wjyy2SPsHMitaMs8bs43qbFvxBp7x+
rO0KtFnqbvPT2HrIn3Rdl6TUrDLwfRPdrwwftW7WJU3QX89hNk6dT/EbVRPZk0HuQhxI6gVgsiLI
SNCtYVTeIDyVOFBlcC4S3qtOw9WD+cjV1uTsujq1tzawGRz2GNUeYpdWRPj0q9giOGqLady2FRnR
07Oeec3rzB0015Qg88u3M+40INC/7TSEYSH8tktyY5+hkq/onYikV4trKMr6UhQhxOvWxWZdVYfL
jbHgm/HfiVUYNtNJAOUHaNo+OAq4j3BHkOhZRCPnK4uxU5CxP0J+Mzwcvsmbq3iNuKeyWf5ngLpL
m0ia04TjEZvVzmi1yoeSgUS59J5pc/SU8ejx5EIK/HyukPiH8Oj0ToCiLlhHNxYDEk8mlM7426jV
kVw2WwtGwEmZA7FYZmfcwFHmreWBMghx1oBjinOy83w8Q6jPXMcTnd1tIYJjsOPBH1pf0L26xwY1
axGerSUfnoStAQYM8ynnDzvoMmHgUQq6syskVBTiASCqKi12AwcTuRyx7p9N5ubPbsQ6N8CwgBUb
SWXtjPRgROach1UCpzotgLo16/TXI7NJrsfQtMoCj4ypobTqktHepjthtIu2MFM4EH7SgvfPlpZc
zW3b11G3TWaR82EjAjfVNDyp0lZvfFn3iQhXfiMe1YGcod3GoXA38l0foJcbNgINjype8Ik63wBv
up2q8nORxHDhBAfLEU0BJbi2sqnNh41RhnQeS20OjaLJzfHY9SxjkLcqZQ8iWIYyEneXrxr2kQpe
NiZ0KGzRbQgFJ5ak7iDVmpP6SLbs9zCNoi2osTS4EH72bkbAEYlFJkGiq44Z56uXKoC6AnZMM/0r
0/uwcwDs+n/Y+DqlVOCHlU/wbi4MtvYu314gztfmk5oUKDAPKzmq4NTJBYOqtUy+/GXo9WE6TdXa
U3TwbVt4FhNh+eqyl8lIkdCfIZQEnLDc01JPcY8dnJvSwJ47mZOF5n8ZXnNoc+XZxVq2waOgpKWM
OKsRLxRyBWoj1dJlMTlIZr3Q9IrEMmXXmxn1TEtx0SIa9OmONp86dLexqL8x8nK8mHQ2VmbncKTP
VXoWtM2z7KkI5RywHFeqhSCDiHcDHSTBB2QcpEp+P750byoFCsGr+ucz3MKDhlgKKyrp5AF3LCYX
J1jyn6apttWlonf4NhkdmP+oJobYkSKPJGNemHDxqs/EpPa+Kdxbbxc09cvowo5GPYzIePGzGTdH
F622tKRAkc/fnTwS2hQsfLdxfJTlCUbMJacvrDDzd33lLoZkFA6EsKBFA4soSNQy4B1Llc0CZf0E
IAznMWVOFYpq79wYrxHDgYqOZa5ir9/XpT3i+8eigKZadsaKtgxOvwLM1oB7yuCpkPYgoYsMtiZO
5WNeaMvdwYoo7hqPU8VP78qFJtZF8aXo64d9uXXGgskLKq06i3yPPQsr0jN4yan+chTzCW8Yk7Lm
no90wpof82Xs105ondIXPbdzMcUX4Muq9HuUZ+3nnESc8FiF9Uddw8O3PkmBIfE/xrkKs1fNzTKE
Q5LflmSPlytpNlAcv1ngtxj5cX+tuL50UUlYk7G8OLN2Xuy6Tl0q7606ZurNfRFLHfAY7k7BO/Kr
wMp1eRbQd3brlNas4V5ZWIDDsj3vHKEpRKeThLyc4zkhcoeNK/dFhfmqa6NswGW/UJnquoui0ug4
1NOmozkJWeMEyQOkCV49qog40GclC2tYsAIhz4bHYR+/HdWRktjfbfNp+PffO/HjnTZGJFnZirLE
4N1yexZIXBw1EsYd3LF4vKQCbpGI02shteI+OOXVxHAM3bPI9wVLmSRTmqdpXNyBvcAovqIOtEgb
04BZcbNJ+SyU1/L0JkiMmNuaNk5+5FEKiv6aEAmSErEh8U4uB2Ip6G/5TnJZFWmEDRWPYkk+pha4
8o5BaMK3i9ERU43nZE4wWPlhi62xFz4fZfR8tSTjrJcnqC02yfBoIqkeQA6BXLiu3UsfjWF6yJwW
6moXwfo05acu+TNO5+3/LOAvJcCYtgs5M4lwmbqpz5GSCT2ECWIk60VoYGbX4YzA5n58o+q93S7m
rkksieFD8LkNSk1dO3tpBqn6Qw1nMgLh5/ROYXmOTQUBczehLCMPPF5kafO+zqIUxuRErkaerYUh
bPijFqOWVEzg+QRwciqpemYbNdgQwRK1phVqJtgcnzmbxudWk25lR8FYVUptn2QYOAqFi2EU1A7X
nWOaWSBUbp9VsZea8JL/Wcvgq2gGwgYBT4ZtqiNiWgnQv/N1RYeASXSa+jdeqZ5hKFNlZYkqD14l
p6x3VjENdLxjdTjl5JazZ8Nt4zV7P5fFueRU9IJQiloxyLr5eMQm3YpTmGxfCt1ozcmzDX4RVc2u
aWYLNsfI1mOjrN1bLun2CoykOIjX9PElSr09ZCUfa6Wsju0H/d/rNHPoSYSTP1gZg/6fIjrb8ES6
5U56mywVO0pM/EF7nil47fZd51YQr/wBTX1192OrZ40dfqTxa/lI0eJaZ4HZ4Wo/3OpkcwwB8gs/
BmV1n83KVushKR+X+DhsLL0FY0KZPuu2+AylCbhGo3OsEmb2/mkNbnHnr+QNWWKmxxiHNhNbH+ML
HxT/ycxS14dMwfR6b1w8pHavMqrIhGUAZkZKHfUAYWZlviLm3O4B9Q6qbmSMQMkXPdfDTveJsRQS
Yc0/Ft7kuz4SOOFXgPVkP7L4ji8BTzDgjMn3Src5nOJHxUmNZ7pi6R2sScksLkXLgl7iOh4fnLzP
E6O4IQRgsl34EckjBek0AMNCgCCgJdOjFp/R0ikASaKPgVUPpqXgafvmh6JscKCKlo2j1+sqP+4N
eySU7xn+eblTbnnmQAAx9dZOsMINy6GTiKKHZtrV5JF40/y+FN3JgymVDMmMbDjMqIqgGsg1PO5f
9Z2s5vLs9L6S5FGMXsra6KwunqqnQr15Ghu+zV45jnDRYoN9nrHJamdviofqtZTPbSnm3d1WORlv
gqreDALrLjzu+IzRx7WkEh9L9kix3dJZ01FxP/Z4xNnp0po5ck+XyU5MD3gzPQGibj9g9usriReJ
1B+wRzt+H1vxW1gedUCZZdgVr6a/nYigxfpd6qer17WG2j6hl365aF2L/Osgc8LZRmlTg2cn15Lo
CGx4E3P9nEB9Cizar6oXa+G4jFijf5JwLq9rCRT3SA1CRBJDo5z0aZdAWb8wZbR0GzC0Y/B+72Bc
WFLnSf1fg40gVc2G3ZxKXs0RPDaXeS+/gBvvQDB/8sQ68z2H4vvevY3C166BdcTokFI9O9YV+2zL
Y8p9T8Eq7nqnAX0QByrdhfsq6hf1kQImfmjAyBOArwpw7iJVhb/iY6gV4doHZ+KfXrpA+NnZVs9s
337gQ+3cOpdO3lgu9GGyDEWcDGg891b42dOp7tSzdVhij5nkUDIr2dWZaex8LoPHJYhAPVQnh/Sr
Y4x10pICly6XM0cmeXSf3TJfKkTJpMVhNcWHhKnh1pWF29LkbiqaMxcx1zyjB75BArSK8AjIZSpI
xFOuUsgmEMgT9upouzqGOyk7/sijFWOceWoAW8ZH3LetSV9t7IHUmII5OCbMVXZDlev8ne6fZ05i
yYXp8vwzXo7V3Lc5H4xyfD/5mMsUc5IFBeYYg1qJ401uV65Ona4RTCHdU8Gke7RWIeoyn257G9by
iFychw4z3xEEfk5ZR13b4Mo6p71gL4z7s7Tb+aU554dd7HaNjVAKC9A4t7U9+qO+ewxLdSqg3XDL
vdhLUmwAx/CYf+KlaaYhwigUeX1isHzRmNQpnWjahfCYFyYXtmomBuXJt51vPgHnrRzQj55fF23G
kfyCMuICUFLmnJKjwHUsLPu1h/Ak6fzyTSrKnwIJRewROy+LJmuPkVXxGF7v2UVH7ufrGY3Y0M43
08oeYLu2TeLpWVKLKQWc23/FxRRY5xGAvDkA7P9tkFBZ8QtS2RsswZ2jRBR/jeq5yxmgq7BI+r96
zMuNpufzZs/c/xvhZfKKzik83dcZKRVZkcoVjg4O+RaSIiAbOZpd/H01ou4v9HX91cmcH0F6Twi4
igue4zN5ZaTynAsVIhAWzq+OhenOHXcdo7gqVPb04VD20xPgIt/LmcSxSrvCRuHgWgahZnXojKg6
GvWiD6owXyEOcbOIGq/DC6eLhU+7HRy15YBHNZwCxmDRX0arNqGX6vicdf+IZAqNsQaZzRQd6vSo
pB5rqx7YWUqYt415eQhEpJS3ajT6glafSsUS2XGKlJNsutoOnMgF/PdAMfVc6FNXcin54/3IxZod
vNI4dUTZEpl0RfCXMXqPqBWM6zqjggnIEBny1Ezj43G/yqqWORBsR2/yMRf6A1KsJJlhx4WuDxQX
ENJrP9fm70pheI6H4lH8wdq+ZRouEpwmWBNYkGxNUcqNjKv7ezXYIsLAlFdxU4ZteI7904OaqiDA
98MterzsD3Uk96YEfwTbDfYs4pA1CORHB+CCGCSxQUdur07pIwFZVkLvTVVfjbAwuQbipHlKJgZM
1xEzBrVZIrT4OAFFOynlwPwkvHThaxKFXucpFZWkqX3uN8eac0fIKMu9OH90LOsMz9+mIZ9WIPzt
b9+l+c7YI2hgq/itsB6T7F00VKEBnuzCw9GPfUKR1c6l7hdCh0JIFV4pQEP0F5NjVdtEjGEvfRf0
buZ365TlnqbBvQ/6FDigX1nMGp0co5RmATriEFSrMRjHsLM8aeofOrtjzTsFRxgx4GVfDNAz0FN4
iETRxTewL/TYQBk8vl7hsQL6qQxzluxc+D3y7j5pXBSGP/d9EiudeGcQDkaCBBxl0qpi9dUBobCw
jhQ5GO6/Mfyqs48Llyi8au5RG55b0RKlpxV7uSdUqaxG0Vk1fJTvgGHA2r7SYURgkhBSJa4vdEva
qpMkdf4kuwt8I6ha2mzgeRKXXSm3LW3W2LVuc++GRQQagZqwHkilIf4pdOyX/dMHZqP0OQBAkXsM
P+CM2Wiu+3SaW6X4aCSdGOis+PVFDrtGVZg85GGoOiwE+Gcpr8l88eg7M+bxijc4jdTQyeKp2k2+
to1DDSqXURS/R7QeCkrahUq4Pw7zBo15OkYqZkhcGwDZFzWyj86z1mAtNkbCHOPvocIzYRLLSUjG
6xXzXiK/QGLMUx0UTfro4ng2tbtJVTm9OX8QbU+flSi+yXqvpBJlq1x6w3U7j85bLNIm4siVOH5P
MaJHR/MMRkjNgRc06heDB1Lph/+6Z//12W10ic8tqF9ABkg8N65nEKzELPtj57gQE7zI60J+1ohK
xGiMulFaHKqG7zfXEH3vq2SzSwRgoEMkiHt8l/ZjDNsEDJgB2R20+7mm4uKXowJxk9AAIKsG6rbt
ftDiUYsj5NKVZbkoUo4Srl5W+DvpnWnu1xKHTxCXf/A6m6J9UI1tywROUH5hvDo7y9Ky10ydOhIH
iHbvqcnvbhdwErL3EuJ6wcKgw/xns0SDxa9o+WY/1EXjjOnGrHRChro1h6qvQO2nwResm/ftxCqf
diOXrn5cIT0lv5mFcidMozEaXEBq05X69I2iLJfHOwuoUfAX4W2lMUFXv0Qqf6XUiDH2yDsfZW4Z
nBLJwLJnoHEnDRe9F/SOPFqJWxlb0joSVceC0diBKLWRb8rgzRe1MUNKYsCqbDfdlHPw8eqKvj4S
ijFZRyWSlLFRVtRm281Fxu69fMNi4uOUmJemK8PgU5zotbSCWLkO0JJo6U5p+un0HHBqD4IDBSlE
a9VMpEeBQAlCr1uhb8gveQz4zv5/428pFzMcGL+cps52VT0Jd4RMWOKKNIobpZdC0ddEUcmviNxE
jMTzOD3sFIMjvV2eaBC8a9W8iMvWy2V1XXYBWz3toEyfbHdCDoRkdv31fEORxVTxuEPQa4P34SVp
Hxd2bOHKRxyxcoUrGyd+KLDoS8Sce/5t6ZV+O4iCfeE7qG5DXTYWikZdPDmAHV9wHIcnshzH+FI1
KSImMpPcQMBGY8JjCctf+v7Y1tpPfNG22CRmcNYdvCVk9xM08MR+Gz6f6KLM6a1wHTNJV9IlMt7S
9rfnkZaZZTKy3eyKNimNKvKkA6nHYxKzrPIZnDh8P2S6jSAJ2FySHalO4eflyL3NK8ZySp9rAf0O
6qxwSjky96WpQWFVcY40D0oAoHtyzugitXNn0ttU6kLMsTOXfwEQur/Jp3P86/axf9w4EZWsAa/i
8ChUFMWQKs5hWO04WsUrv3selORe6Eud3IL3wWCIZnFonjbvNK4VNCDY8D0TNZExHbXew/HKYlRx
yyCQf1FVZquCOLwE1mJUznNgQi+nZzQYtYib6FyfP3igzuuEM8J//CpX6eFkmfzgqqXZgS76Pj9T
6pvlKh6WNupNhOnXmaCo5GmFS4qWDkJJzXa9PWtE/bnRgP7dG7YFS1Krf6o3I9LIjcXg5PvAl2pL
u4sznGCiJ7sUkwypH9utLtdT1l5W+AGQuETl5OE23d5iWsQLfxt0DoBWiC5/VlPsFz3EdlaGnz/P
Nco3Xnhv6lwn2Y59VX+AKvpisark1USoSA5BvvuhY3AWvD+is8twCZXkSBxk+VEsEWce+dTOdmH+
WgW2WVYezn7VIPOHUZioNPUYmvWKdOCfhWV+D52LAFDa12iuWYQSq2Ri2RjBd7qbHik3XIN0cBfG
H0YT/W9vUZqX6qa5Kg1r0t2IvJEqsdTqBfV//qHR/GD/vvCsCpwsc7x18pUjG+0gS8fRdWJLHKAw
pQxAUcJnjOkjGA2KNmnNwjzvx2HP0DVsVdGXEpILUDihMsPd3CFSd7VKet1+p7q7HXvRmsotgC5U
wgY9KKavq45n5hk1yCDSmuGSms9KtAuz3jBEF3i//4ZRXN4yzZVigYefxPoNWm6BWCel+JYEWtK2
ChsiptKLlxbPlszTx8i9264tWHZ2Ay/fU1u8jVsBplSFWkzGSBPwUmjtoI8EyuIEAkDyxHQ5uUlw
RZCY6Mw/FDB1xehDXNZiI6oGckcxgN5ULnSMkxS22Qoze2n2mMlNdmQOP8T722GWfZgirH23MpyS
31PLuj6zWdx+t2ontpPjThwJzv8Gs7gkHJkIgUt5eSohvo8sEb4uG2wPil/vI8ZiSdjI068BARen
/ZHSDKDj6eWAY6m1TcZpaJWP0x0S7xs7IRQkmaw3uP5HPRnG4np6DPTP7eiJEHu3h2cPCEaoXUWW
F87GFrt8QEGhOju7UJbO/CO8DdhfhhKmCpbGWCFZISAjdgyeX+ds50qIh7yEuugy50J8U+JBAHgG
MLuJr5b3p7pnQ89Xu3fGSISYe8JLy3T41HGJYiw9g9TkBs3SNw17k52vh9TQNBqF4aEFe8smaWVl
RAvsY46iClqP3bA39Yg7xKdgTo2k8dyfVIaKJ1NSeFLCGPje6I6OFfZFLLnYcKR7NhyBjs5r2otr
Y1xBQpYb/eWuEdWteBKxMM+mBadBcB+/NGGrASdYGA1VSTHZHq5702lXqSkuWyKP+B8UNBwQQVwu
adER3C8dKPfJSbQ6dBCbEEXTpp3NthF9whsm3NwhjT+qspTFabMi8AzHwAZVKV9I2klNvhNPIkrj
zOijS2Ah+iFetLVknbOqXc7j299vTKK3OVgtyZeM4IqfCt4XJ4PVSCB+Ds6hCGHsKuGqINJ+wH9H
tcY1xymFjFBxEFkkoCLXqYZSAznp2xQCQRWPT+usqHn9kClWGOoqtBBDMjONPLjDMB4FjdP7HGYH
ZBiuQXt9nWUAfW43nDLZArONrSHseEedNhwiu1bBJQN56WnC0VPmgkAwNNjh/78mIdQmMD6uCgdz
Q8Udul/vqxcZdfXprKqd45hdijpJPGWvkBoWgRyZpcWpTfEIxEpWE3vUJBl8dDJ+enCwejTglF7P
1719HeGF14dp1t3jq4xoYE2va0nw9ri/2qO3n6HM30boKZy7meuh2RbGCzbReNctp5KJckzqu10g
mw0xgv81hxPUDKe/oa74HesG6BcvZwz8GieYLzE3+fNy/+ZXcOMBcPZ7i/d+88W0bxgQ5uyf9EjE
PvfAhtOXE5dh6HjAC7UzZnUn/xhgA8l73D4VppgvmnyH/lRHvc0pJFWWflWv1h+ySa7Yxx9GNoFd
0QW6x08IPb1W15+LmW0W7BhAVvTKOb70jXI39xceT3HVK/vUu2jgl3lgOZF8ZGUM6KHXkbKpB4o3
f6mh+NecZ6DiApOIuyGM0LcYcvzSByZUUJA6ehWcT0zTe8FjjJvACl627U2OMohx8lv2qI6oWaaW
HDjYhxlwoLjX+yZcj80wXn4BzRJmYj+/SOx91LNuu+tuz9pz6UNcTiOoKa/u1tWKc0bKJJ+BgWXk
fky4ZjvjePAJVNAJVjrmg1hyFb6qSIO69x9gTu3i0g2ByI7+dYC7prOw4LvSCPFdw2A5u+XVZPJe
oVOkbWOJFEDPkoozBdjiTZeeAfLyLBjjhsr4PM8B41VEPIGEBCWc1QiL+WAAzlDnKyGUSER+QIVP
coeF/q5GRLZfSZghpx/xxF9mLbjKwUbedrjtKI1OOJ2FwKckiPaotVQP6DO+zf0Mqsuz0Q4Gm4//
/yrdY+vHkvuHf7N0/q0OC6X4zzq+5XdolLMYL+wNks8nVu07kkliI+a9xe1bTD9jZBCXjopu8Bf8
dj6JBPj+QvjHSbR7GFB8I7iCExAlP9f7CwFbita97bTB42R2C8QyjnZmm+5zB4ezm/l8cou3UQir
8y3WHpP/tx+BtW0k7KG0tXkefJaTI/z7nmSjD625qaaeyOSmixK2j4Z/K4VWaXrR4ZS2B1i0VKoE
KtwzmbXA5vRjMhuquTFhwGoM/jHG/SUFcmMezzPLKiWTLIYEAkBWPqatAA+0Pj5uZCRw8JI4WOB3
MK6W3g4tiYEKZIyL0OyNsEM0QdHzAvch/Eq5WsT3q3beTjCuEIcqckj3m8yqizcAtci6wZsCD6IZ
YMPlNU3gakUmeHvuHNaSqYXT8cU/Pl/PE51JyYE3Dmj7Vw1lE8rxqlKTLokO/+u2xCYXEpy5CEBc
H4dTLLGwxZopRd338t7wQjlale+u+MduPK9lDgA7/4pRp5aozjrjEJjahBt2X/Hb6eJ1qvEyZg3n
r8vZbDUcWU0zcSoLrapHMcqPphOCuEnmgs0z5XzGZBMsCaBU2lLnhRWAdF6u3DvWjtPqIZXRLSiU
E3JFVwYA5phDelN7ir8zVKJyOt7DrgausGok3mxeMVGaBxBb7lhO6fq2LrAfszSX2EvS8VNtvypY
nHA69oO7H8B2quPTF/PDInPo+1J/hqBErt/DplwQvxNIL+JbhW9aMvdogf4GG8GZPo/ujRlTYSnT
grcPIZqseNn0TLffXIfPhLE5R3XN1psKHT4ptmril5qR1MfEUjHb1kwWIijR4IOUwxLq3Kfw9PkH
f6ARNMutWdzohtXbvYO6NKto6MkxH2oQAkCGvAPs+El/W/zpoCXZJsmZAnGT5f51DotBbDBMDhLf
x0J4X1eO1MZff18GrX0KuifdQg0eIZNPDFtdW9o8YCjuv8/0CFs9UNAzHy2ylzXFbl7UZvPJ8liy
kBcHch7XG+JJgQ0hEFC6d8qWot8TyuT7U6U6SZeTxJiXVolCPFvx3ZAF7oA6/SfmjffAGucX5YbL
gxpuqgTnlZY0DNzaT/zjqyf2nyrEJeH4yOv6mDJAB6DwXtGCZ0dNVnXyNfXJYQVUMX2KpJ0tT6qe
LXyFTOV2eBYjLdliGT9tUAADOX+raKUqNmQsnnhUb9iPSs3rbWmiq0M86QvGFGE+k2HuZ1upMGq6
O39v5AVm78Cj0EXbJjiOXqI1DSgCzaLmhjleQVDiPNoUAFu8G34eG+EPaLjnW1/y5n7/l2PW5N1D
IqGtq8BUn407Wd2FStJM+TAVr79LKftSKDrop85TmGC5suT3PlyMSRvmrVjB5vDurLKIY9HkziOj
CQVnl94X5emHBETktRy+nFTV9R+swq0LFFvSZrdeZgtbS9XtrFDYZsAIQgDiX7OX2LyOTRQz1t2K
xokQaxDV+FXCgXE+wap9eS/moGzTFkBKhdktosnMhAoAW1MqGBNjgS4AbZdldA8c2miSe8exgRgE
qoCfSJq01MhE8B/zLCRVd5SUrNt0YEcvSKsFpuYMiBjUOwHkI4yuahgCnXw69TgrPhJC35QCIdmG
FC/TCo42mA8TQ5gkVJOpXHsRV8/LWRWtB3oXrhKnxP3SWBX6IOCl2anRVDgAo0CAi6PaKbFJ+G16
HQGS9xas8skbQ8bxtZm4QScIdN8BSsT3iLzZjDhP0GvPhmMERuvcuk+Fs7L3ksH3bbQGHlGpxKXt
6NgP6UJW0OX1un//lwGOl/DhuFCoxtMYSpvgYTtGg9sbn32SdaFRxwyIwL/2JiGcpmu/oPSnDZt8
7S0aV+t9KmclDPwnavswsSn/tkskGX1SeQotrPS41QNi0MpRBCC63H58W83bK9jNw+BMPrr8NLpI
pWBzUGUM4IbCHPVowtn0wsWwEV7S9jKrH4VpPX+IIuz92tUgBZMMfIdHB8t3eupr3uo/YpKs7G1y
G4TvZbtEwS0e9CVAP79CD13I2AlqkFdjHfCMSXbFhbUiZ9fTdbEp5lc/osQtDs43R+yzY4pJlhpQ
lSOL8Zz/r8FmcuuL9rC9EOzMLzfkBWr5AmKqaWM6+WohjfzISrGb/3Qs3HNGh+ACUz7QlGBgy+Ff
miTQZ3rkKzM6rC+eVYdlwXACWn20J0VX1DafMVYZtl4PBQQfOZxYDXGd1HvNnknNLYknT+Z9oklV
gQ5xsx6OwrU4lWlns8VHqnwsLlHepS45oO3fCepJKXpyMHT2Gvf0DQy1Rp6ELpJuhoWhQg2MdSSV
H0Mm+z3hOFQ669ov7FCi5Mq0rNKXO0CONEFpfuMVkzteO0uaMBe4pX+SC9fJVTXB8fcFDO56WitO
zt0C5kpFR5BZ51bfSBybwgOeoM/ssm0k70poci/jZ1niAeCpPyPcx4e3ktCVCRLQegnHlZPBoPWd
7PciMuPMU6TeW0ciQlH6BLfW+WnTDjVzJlWzmSbvyhRAfiuGh7lTS4Lhl6uHnDuptvM0N5fumpJ8
1CK2W86t21pGa0mFNsGf/YU5ab28p4Y6pQpw50T1OuBM1RwJNWYpusfWjkEv5S5HY/vMGFXHtYZy
5ajN9IyRC8Ptqsep6gqIPjETOCNGirpjKRRmt244xyxkB9r1BHrj8zLpslYf3m5es6EoI713Ol2S
9ZtAd+7y8ep/f94N0Wa2gT3GYrB7C49rvCK1JSWRI9Qws14UnaAWtJg6vi0FM9z27lFKaMkPklze
zh86knJvy1GtmwHoa89J6SlC+nKsbpPzeMZ3O+nxeaMwNatk8cZpDfeNoDfljiBlaEXOTHWDoefc
TgQBiwLs9XtvxU34q52Oi43vs911xTMS6C7UFgrgsRNJcZtcAtRA2hrQj/T8vbkX0E13fzwH7T7f
/OtZg/lX/RmWo5A9hjniwGAxzSZr1bEY5Sq4NwIpXVo7Ynsh/HCT40e/hmM5CWame+BwK1bYF6oL
FH6TqJEiVTn6YR2bCcuwJwRmqUv4jQ3lAnGJHYi9z4dIsqDWK7yBcIUvYU2hjZq0sBmNBsynN1LX
tBPguNjnpbbvM/4Zjzrrpully4PoyLtVUaTXc+80ZMA4xCTk4i8rWpDSt8HRbx10+qgCyjyQ0jjd
Gho5Xgk/yQyKJ9WtZvzMb+ieLzPsSVJY+35BsvM2GUsLvbpMf4Q/R9a08FZKmBPAvtVzSYnFDtzZ
NP9PFEB11AWWYOa2flXZllusjrHQzTtUjlN7d961EqHAQc7q2zFNWDrSWWi/wLoHlKPCoCcVSrtq
OlaX9Aerts+9+RpaBCwIyLrLwBiSz4pGaELOffozyLO8sxI8KyG0nqoJLZRJz5EkVvPGd4IY0PRw
06EkQIFLihMu6JYsAHriVv4DeCRt8rnZbyVqe7xI5+5vAxRTDHyY7Lxfh6hPHXnrD1HNspaxkGfM
uUpXWe+7sHyy5bSyc8JXOzM7QNkZAmy/OKgUOavK3zxpcDzxZ+IXITUK4mX5ufECLDsN6oNi0LqY
wMd8qwG2615vJPhKoysy49J8xRTBgtVaESyWozqGZrctD+NZZIQBuuf7yhfI3cM2juhDTD6Wt34V
vuHSMlNGDQlGmXkpPER3ISXQUaIT8GjnOdtmcuSAeED3WXLyDtbOdgdmJ8Dx1ElaiUBObPUj5qzD
JxzxqSIRc2leRqXNNMGiQRlveUg76CBkSAq1WRi93d20+xrxGiuB4zOMVIbv4q875pHLvaAuHxbk
6apF/enavJes87LKv91UzfAJTLDv82dZnotDZuiVJ4ofB2tGlBhLz1dIgSGCG2dRemjWZeV3jxll
1WOHpqXoYThN/cdyPDxGEJnpSom6iMKX0tNLJYZ2SnjYk1MUFXGvfcT34zArOTn540TcuWCYQwIa
DceA0JALRQdx8O8B+SGo1hYfKmvDDy9lImu8YqDFYmt9+RoTrMv3JcAWhbE0QNWbCxm414d/NC8k
kUhgd3DbHs+IUbs6gTnkOAiUYP/m+s/heT+jaGw00eNDedKKpYfjtIF2sako8CmfBMTdXf5bWxuV
/ib3NLoEKexcssOyd5Y7uL145qbi/m/AqyHCfmpKlxqz3YMt9/9mGrf3DJf+TzuXhvIzABy18op3
3gOKmxL8W+1wEhe5h0E9F1kQupYWHOc4n3B3Joq51LMeu3F2aCYxpMWiV/9pJXsf0xvyj3EqI7ht
ePG+sQaYEDaAM6qx0jH6w5YweaSRobzjy40Yh2QLkDX4jqEdP6isatZp1VMi1em0WUEe1OjR2GXB
jntwqD7ZqZhpcEWI1kMtEwkLrMejbz0sz7CuvHNyd/PaSfiOAWxEPXnYE27wjMeds3T7Lz9M5din
eQ/M95eU9ICmZKQeF5lJL/xn91Xq7ZhRejN5BXVAHnrgDnK7diWjMiXN7bjgwdyA5vIAIYwotSPA
YdakXgIplvxCKIwpDcIC2qcGu6otMlZdkNy9+A/kqhnUc9w77e32F04BlYRlpaup8WSTAwj9wov0
NZaGM3VPHpEwsK0ZV5G//Vm7FjJH3H3G+UIgVNE+SFP+j4zszkeqwxE7XM7TIFYf8ipBnQTMX7fi
lsqZwtxfmKyV+2jrCuinmGCtWVQseKLBcOggHyCY2n/NsH6NgT2GGYRWdzr+DsAY0ogtbvJ2Et2i
AA07rh1fgbItIYe0I04hlXVpYNAeDsJex9wZ/phpnhyRjOEE3nenGv800ILDqRp6szq477TCX0Tx
JAGaTiVJnvsE5kuUrKAV48P2XlkSV8kzfTpbSvYSG2Ij9AAQSAv8rY5wdGXf1ELlXgta7f6exoFR
Nq5Qf/8SG+qqE3omPojvY5jg+7wBcYOfUijik8yPG999IR0GElXByvTiskewovKcG0KIRkvSEYt2
dLFMh0xD74EUcqBrQkcXv2luIXduGMqX6chZvbCbEh6JSjCTLRBNMm6cJbP6EQdWZiCeCJn2pNwc
MSIMsvsmckrDZaZeiZkTwyNLzPMdWQ8M02z7HLKRUXcjRO1wxQZnulAKgbv/K6Prgm6pHuZPdoAY
LvECrQSu0jSCYL3UVosyAPo3/+J8vuQtqey5G706jKu4Y+yA+Bp2mkzhTCEQIVs8flv7EtHq7oks
c2JEqw9f7cJr91Wo177/DUP+EQxx2k5Q+IBpa2Z9xQxymh7QvzxYxQ46ShOR2g4MPRM8km3ug3GB
TsXhN+ZuW+wQ+sHYFQ1vCc9AP6icrvYddoVol37kKV3/Wnfe1VmLjsi1eM4lSLegmRcJeGONVTgd
YWt3ya1s3OkJCvaJOuyCrqojSTjxLAJ2lrkI7CVEXXyQ6TMAqhNqJQCw6y7Rx1ujrNNGCjZuQx9e
/52lpqqjl8DJliGX5mYcDt4I9bBbZdd3/5zWWRvbA5liWRdRQ+OQ7s5v5ZgtpF5GZSFQW4guxCVk
4jUxy9TNLh3D5cK87UznKU5jqmhIeB+RnMnAQtyTIz2uv3wUo2C3GZ+BJeJkiV4J3CaqrTKwl6eq
0KcoCrGOcewfDHTjAd3TmDFzdjwUclC3iKofZj953DYuAJ2PwulmDBTRg4/nxFk7iBVATUgHSeCE
nh+jVYmddFiSpV+otaBZN20SGhc3VzlgBPhw69JicIJem7zz0ylqNSIGu0BSYuaZ0ECkwbaf0l+O
FE0a0SnSHegdr0i5tbRebjLxik0FuuWekzYW1vyWaJvBk/VPBvpxQaht/lwRKKpfSBV+rjjhN82Z
ArG/Jyftf/nKaHXB9PinlK6nZFfk+KY48STCBK9qhhIqDnUl1ThqVYwmMcj0+7kyej9LaYRhNaBZ
4sYa2ASdNxhNGXvUfIPAuAdnLbL/Wfp/nxbqjhqKzcTFLdUwOujoKBdpzVMjZJUTy07fAb1jigJH
quct2JIy6aTr8znGzwbrr6Maq5JqmPwP0x5Leur7+VfSJMafjd/vWu3FCDcEaarRwoJr1qSOK7ho
lE/7cKL6vB3XINl2QJuMG5kyxVwv7FpITQmKZB+Z74ohKZBy4vWOrVsQv8O5ADORZIcx4JlU2iOH
pb3CJqgiHkSnntMorJO906R4QeldDCXVNr8BfBNWXCwv0Etbu1OBjngsf+UVHGIL0+yLXM43eZCU
8Ig2QFZo/3j+JqKqXOKo2Zp+2J7R3ikivbaq/PMF9NoecqWPej9p170FWuKOH+4kl+2XlnLAtwMv
cQyT5eeG03MtmGsuajbEHRMsSCAMDxtgsF29zV7SCcJRa8ApuCHdyDgmxZqZDyTLOkGoHmo+Lg8c
Ps/YAkkaXQZ19dvz0QoXhoUn3sCQRd81eDahc/zPck6u81CGrm0MFuQCSTYDr8kpPWJpLzWAOL0C
Cf+kHV0SmZ9Exx1gAW+dEoQV/e7LE8XOD5NaBCxnWdUdAF5SU3SQZneQ5yAsAtzz0EibNJ7NMF9v
QIyFftQrToCLX/IkX/37nd0DQZn/NfB0TwTsyhp53dyfjMfUhe/hSUimuq30iNJP9sQCrIR9sQ+y
PfNJU8lii51OTvIltEVpOaso9MgKC1xyAJk9NFcKWIvu9bTC6N2c2y5bpy5XogdwYuFAKqVxAH/i
4AxaWX0EIme4FBx1ghbhy3nFySp9wNTdjFL+ogS+AMjRAZLX8BB675WzOI9SW/FtDrWwH0e86qkB
YhkzDhveJZVDwBEh9FzblfjJEp6CKOo63kShv8seWR0vS6N0Ff2/CdLsMn15mMBsOjXgtCqGX1bh
U+W/7+W3M+cDecbRyMMnhXwPAWSb0W3iadTzzwZ59Un6N+ao6acZ7gj0YH8yTabJc4LNgFyS3cZK
ZqSr8Vqd2Rv1DkzRPEb5Sf2rWHPFxtJQLsPG6SWuSD3fOv7hcf4F77Zg3UiDeNBijjtwpoVjeZGs
uQOAKFy6EiC2rr85EBbIeQSYFYDIBx9mwGZYWqLNQ9oJ5yQARSPhtPsNk1EgzcFUIbVSUXJUsPHD
vRREBIrd/tQq1GoS9IEIqDIO4fUER38QsSeoYy0JsYfpKu3voUA1J23UbHFjZoXk9F439xS1TmIU
u9YhIKKE9kCRzYFRMYZc9khdjyEyDbWTi/C6RJeCiVy6RPNaMCEBsR8QZeNyx9HylrRGB2MrK6aB
+gy9UfeiKZp1HaUZjOOoZNt198DMRY7yYAZmUdAQN/JTQZwBt+YWEWKtuzV74E5iHut1dgyy1CsJ
zQNSQdjg1PE3fClWrpcER+rsFzbnrdttgKm+XWuiSjHHY6VUzFXYdIGIN6j9TmwB79qGvjz9occl
Iz1CdFVLr8gQXQtw/lPcYG5lLqNvW+/NF+eZkc+WV3rm3WILJ1joTvpIbPuLkA5KdYaFwdjOYfRB
QQkPLV6m/A2YtfzMa1BjaovnZbhTXAsJVjnNE3L81CrAx/wZK2euXBQrnyPQ26wZM3Kq/NJGbaqq
YlGGEhcKi2M608dDfYyHagvhsdUhXM4aGOBsec0znjE33iHgSPqRDyTRmeImo/LGc9RUL/US5ZiS
+VmRgK64I2JyK6UIt1PalURspP6gLfWDcprMXLI4BgBagaMf8PNre1E6RDums5QYfAZ2KN0wx0kI
TRZJ8NCVMICxylrms9PN8IgK6pTgp7FGv+JXUlX75TjiMflaSbN8WhWsN7uI0nhim/mhdzm79ysI
pbvyKqPlM9I3SV7nVJrLhpr6wG/YpM+C7Tuvo6mh+2yjnqFSzaTQBIWXchiV28w88XuLkPAPVfFQ
8gOc/k35blKOc3bcrZRLzAnXT6hjBl/IrwkROR1RUqbuE8OiLB3Od9lKkjMB1348SyML1slLUlf8
EbwUhvNmAstENzmI8YwIxslBD5V39T32UuQSQvNql768yR/8rN+aQ38k9rNfc5ntCgyUsS1VZ+cN
VlLVpg5m3X7qzYv8NRCIjaxxs+t6wSGBw6/XpPt+yvIVY/Z9dU9i/EWfT5CnnDQ6pkWt209jZGhO
z2cwZBGGlhPelH1EFcU88HlQrhepviFj1jZaa6epIFKVM1t3tnGleACDcCJp6wORP/Zq4S+hwMWL
tCibCgLxUek7rHz6G4aOVJjuZXkTByRlbxE4oXOZJ0+60DdG2k790RArkMHERysaF03bCOtFceTY
yvjpz9DmDwZAlmDAu6h3IwwWjiZew7lOn5Nzo+ca2jJ46GKBe8n+ozRZX+YgQtgLPau2zIJLJG02
Dx5677HPGcgXo7G85kG8XMaWEDVtDDKSU+4D6WYZm1OhzDoIvZWYBxHrCXyMoXsgNOHfG4Yz3M9V
N7HkIq3NlGCsrBSd/ZYBBhJ4W2M/9zVd7ym3Vr1+ocLIeqk5spb6XhSC4U/7/hn4YijFsqlaxtq6
FotLEX/mX2Ajqs44quBcw5GWHoxQvfa3D6ZPjnm2+d+OghcqheynodegSDh6ahImgCapGmOyEK0G
o4dP7HlzdQMm0P6z7TJxyEK5hLy96LybDnZY2aWXxeerdEGM/LUb0ZtXbzUuEyzXe+vAqZFj3fCz
OFF0pQtYhvuzHsfGOKgg8CrKASjtqQTo8ZdcpJeDomi2ANSFHj9GiKABOjsfjTwFBR87qJyt+xdg
v06fSn1ctLyT9iD3C8Arxrf1Kn+9ua68fyD016Qw4u/QfQwM8oMYYnaDw4Kt1O+3Lc2QZGpHj2tV
NeO8TGJyR4De8tS8BSJkYN40+55g8soyF8MeLkdTh5dmYty6rgTATSdovZdlVy/jGCW+CeTV9ZQl
2x7CznSJEenpvuvGXYVb/bm5PRLCfik23AlyNc7e//sB7hJhQrqciPtP0AXmmym2JkWSLS0OItj9
cIUZwC0tx6Ne3CUy+uNlM7oXnh3Rmulz1kNHz8q5+jdEpcHfr6tRlq8B7rB8KMAQyqcYBdauVRoX
vKF5XhXkVrb7XBRsEMZD3ZKKFA8+JJlvg/1af7uU10FCjFqAaqyQMlaUWq2tB5O1KntVKwc2SYml
AjSB/27wSk2Brxhln3rQTotnqoa3YZGHs64S6I8q9zS6flwHXx1KUdYqjQotjjr3Y0zUKX5JTCnM
uMxTECdPxu2BkkwJhw8GOhElDxjOZ8AcL6yxiuHBGjIn06oaBNW/4Om962hzE6EFHOIVfDJJ/FAn
7CXpmcqQW2Ts501yTqJozurcROoLM3aZarQh25HNKB+0es5rc49/s0aLNqBD9Sfrh3NQDlP+676K
X+zsrBJoDy9l5WsC6N7PTrkt4lQVk7HJBOOPtVOnTiaB8NRiuWUVNJ/DB/uYHGCcs4mzuf1mcxnB
fMkRbAhE8NHFcfc83gA5lN1JnnylyUGE1IydGJLRP8A2dx2gfkAYn2TI2RPHUzSCisY2saqN1k6m
ULrhCZ5UkR1FJYHi+ajr+SnJUGQGSQjYBLRX5RXRQYvBHl7qR80K8oZScDXVocmP9seT02pRnTZ8
/S9kNzqbbJB/4JmOwLUWmR4iVSd1JIBQT1410wBwpM+ZtKPJkuOul1R2YUcQHA9bjNJ7I8uuRIAN
feqFZbWmDouM2kwPOpBSPZdSv47L3DFcr0YJeG0rdWggNHr3drRuQAT01K9IUN4+Cnwnh3SGkI3v
/FMzS+RhlF4q9X1dplveHKRJ7yAWZ21PZkrcfTrgixw6dJUrRPjeAx+jifUR3UkeaVTRR3E1BDQ5
xI6c+HBnayRO1/DkCnZ0U35kLNCmUcmaovGp35Dk1kfp4PtPkGAYl6X6eofC5DYF1r/VPQI/YIHX
YkesjcygTl57tVSzjq4bFnQW2oN2bzf7B4/6ftMyMSAmIsfq7bHYh6V/1dxLzv8N7jlp+7tc439o
nqTrm653LK+2lmDnSxF9EVwnCATOnU50BT1B0Eq7ab32fMYF30fYFLuTJ7lb5qwIcMymGqbg3KDO
sSywHHUGXyPyNK/1VERErl5lF7/U4iQWHAzkDqFUTNwOhbVeC853ykgnFw5LRf524owlmuY/RDio
agfQr6I8dQ3tj0wyXO9Y+NCkPq3rSnvUugnUN3FXKsTWdyFEQyyqXosY3j4w7z4MTAPMrsCzkBhH
o0HugaEN+3tBvKawGXikc+fn9RZKlrdjG5iqg2/+IYGlOK34YyC3CjfmNdoOPtCxWndUUat5kD8j
YuqRnUiIHEWRpRYIA3uKHrVGUYpe4dElCiGRh8FyxA8PhXBINsYaxFs7AMXHEgRtHtAqHSiVlgu9
srj+GJpO04wBhVUvnm6ZdOEl6NwV0EYpM9j+DSWO/nyPxsB5DBM/z78z7w8xIGZsuGQvKIz5e7j5
T0eioSlrqQYIL6OpwsEzif+nv+A6XWHaf35AR8DrBX3apT4BDMb+qf3J1dLC6Y8PwwiyMjthrFlZ
yMxo9p0BbkPpTuTk2eM4P9xk6sqStskHx2GKV/xN0RpU7ahzZWFopAfDHgLl2KPO9QCtGWuSYaS+
PnfT6xVP65DSZe+NjCd8j9sEL4zM0uEiVq6KyMetxeEr7FFkusSxpe9amErtB/qhqfwKT1yMKZ6P
Wy3m/ZObQ1eNzygUL+Wb/Jx28LNnF6WjKaSfn2Beg271nIZlfyi9NM23VOCHWY4MoRfyZ8WvPrdx
J3cNQDvITRRUqqo5ddrnJXd/gMJvkVDuqpV1Fdniee52pvyU7tFnpJqn6V65mn2WJgG1+EVQ9ESi
f5GC6HD3MEQ6wjCRA+0pSJISmtIOQIvji+B5Fpx1rvF0G1gN7P/B3aEDa3a/BDnhIz8pV7A7X33B
N1ziZGfTTQnn1S3Z56ArQDKFpyLkbNxyIFzp669/Q2ScCAhdoBpJYOne9ArJKZ3q+us1QHbdXFd9
1eKRPsoUfWufQ6wbvhNyOxVcvfA+mK0PDrvo0EC26SF09hQhKICiKMaI4hsylgD3QB7jV8UeI3u8
+Es1Shgy4tKOWyCUPqTB6uM0fbRXtijfbRhluUPCPHvkUxm0Fywa8xAF5m8becbtCMT9isZENlzD
b6AiyLWU0hWZYq4ebPO1w7mhdfv8SP32uAwwNlB9nqGyZ3QPhmL8XVHfcE9wV1hvo1rbzoaSlA/R
EXXMStnpBS/yKQXTyqyITGy7Je0HdU+tdKRIvoGUtltzge2hTuXkSIPCsrUhTqLGGHmjfesv8lRV
jkE8mXPbVKlVd8kF18aAk5RmpUfv9QN1yrVYjnUX16bste4sq+S41LigYjd2LOW0NzCEIpGvLq74
9Ufbu7Vc+PFfI3z0E8Sn/3ZarGmdSmpC1wbWrKt6FWvAALIuDR9tnlQSP/LZpI2NCDzbtXLKzl6/
tOmJOhZDTGUeZ2u+VMn8vx9NF+sJiGmCNUjwZ3WaWVZPmDMbHX3TyIMx4duUtErEPNTVLSJZwoQb
+yh6lKoHNA7MH8KV9CnUr9iUt0hxBiiWbEwYGSIMlF/Lxso0rF40CLgFkDELLA+2IQnjDjHSClCd
XUYTVU6EdupMw3y5c2lqRNUdhQ4BIxbXOhkEqb/n5asN43NmkUz6lr4lD2OKkAVfwYQ+amuOZ5uu
W2fZq3aimGezNSW7v1iaQmAo0BrATKkUyVyZY+eWDGD52Br3NBmC9dMb1FnlxZtlmZj29rZnassn
bi6zM3040OwMFzB4aExSRYiUqmZFds3pO+LviPZmcESNLAPUOhu0Y4NgspA1niAQVpF1irS/sPyU
om8mNJHN1zGhG4zZfM2XcCRompxsjqHhFw41/DjApCGXbJkfqfiOM6JQpsfsNwaahBmXt/77QPwS
wkT8mxq9BVg2vXhyaPIffgA6sbXwYhLQKGToenv1T6Xkrmam4pT7Y2wtxfix0TJr9jGJjKaaHsgp
MnZeONiSAJE+Iy1cUksJSFEh6EAVAPa515SYPogcz0IgdUoHF7SoKrII6uPJaAtsAFQsUw/B+qzj
xWgLn6QT6XYAqEFd6b8b1GSrb1UxXP90g0slgyc2arGtYEfZO9gSt0Wptz2wXJgSc9paOrHwG/38
Ha7uUyUMCAoSAp0BxeBhKW2xv79b4GmCpOew6bHj7umK+v9priYQZNxffV7di0ighBjKx+7MHCW7
9luN11FxOB51cRaVj2fRKFQe699r5zIRWUI4hDaR5VgfY+3tkI1AtDKSGCsgfrrL0cSoR/AHVyDg
GsK/lD1o9Yn8dMJsCp44u+vvN1S5X3vElHGg2MM4BQccO94UpVqzy2sD7YZ0cLg70yh4qKpFvj14
GRZOPrxWmiXzRqBFL8psOFEv5/aoqW4sBMkb/lwg2hcwXy1zwuUEw72k9JiKq64q0eJYEcxau7EJ
Gz3MC1u53J9FrUkZNWKC9RK6QXDyhsSz+W+G6edIXj1Ocxd3qO9l1wnZ++9LZUM8NNUEuD0MLdk0
d46FpKm7t93dmD7s2yBb61RxjotcCUTtC+1fb3ih99z/yWB3HWN1B3UfUJTY3UjzXwbJDLe+SKYt
S8prBy/qBlZtW5YeHuUjolmFJFvsvTHb0uMJ4ye5JOddoLTFtAj3R+AUCJjLTuXvG1dY5AXN2Nky
FVh8yl5GP45YIY42aQV4dKPivyM/34SU7oy03cPG+ABls+a/SggkpH9Oaw6dpFgs/Y2ukPcoTfoB
29gfoT7MRzBxHuphMA26UE/Roy0r2+0s/+3UWoi/8WtGgbFvMk0G5Cd1NzP+gMaVfi4kVJY3fJEu
f0HNSYAOEB61zWVIvtzwfTZMEU3YQH58jEJ96BbEsssHs/YBnZzgpBB7pzgBEFaSht4ZTaWU0L8K
Q6J3oiEfBFB4gm3aPUdmR94ZAd16LcIgnDXOGjOK3OQ2dMRAUhW4KGebfH7o/lloqhItwkhzpBuP
+PQKhkqbS3nR91gUxZC5iw8lOVyZDkssPL6s4E4EGNCrqGuvvCal3PDbhJU3mxadZFW1S76KAByO
efG43ZO9OKzpkvEU2XQ2WhmTKJU434u5JdDwWEgTSjhG2baYHnOVPn1wa6EGXj/JZ6rN5Wc+C/0p
ecojTaca8NUEYbXc0BhDOdSwyT9brLPr076AalxGPAxxQeaARfjIlA+3HLfY6FJjlITOx1KXLmOb
Wf3VnUC8z/FJeN+5+g6Jn7kSeWuMHj3/fLQhxT1gKbH56y6BoZfS2lRXymtsxnSpDfmew33FI5Ro
HrUiQuA8ym0R8B8S6NzktV7HK3zcShe96xOX+vRjxl9cmTjUudiFXQf/dy2dow7TWnFcPLm512C/
BrAi3eoY4eJV4xhGadKCFIr0++VNHYJYDd25zyOhIxMX75jnw5Anx+ja7e+WUcF5wBPc3df/Njtv
mnegPaWgDSDVyOfiBXzl9eudPezDpj7pEohgi4U4SvzMq0cXNruyIygye6VVZ+eJGSpebaTcR9Wy
OJ786J1zPGk3SRyzLKfiMPDvgzfuUC1qcy4t6k3qYN090EjqxrDXyl00QGvKEn7AydH6f5jOpYfc
mI+HvSYSjZUguP9pNBju5EVhnu6mX/q4QCh6l3GKaRfFu6ddxIIVF9e6df6XPLNlzu6Cc6k4LUgj
1Hs+2XSqWRi5Fll5eDjxNR5xVTwKTQ4v2yXKUe0+544LpKV57XSd9tuk3PY2DFlmeqR5GRAfGGLj
1F+uVaNY6K7StBSFBwKN3OZNcBz8xasEzBvJ7pUjl0zfOYh6ICOQVuxnHvIyG/pjmnN9X2hB9vq/
GJIJv36cpBlTjTBMj5OJYW5B+Mutt5la5jCPwaq6ayiXiyivRsjk2UtumHQ0TF2dU5uVeiXk6m4o
aeCqT6M4SHApvVX/cCVGDIHGlYuPSZWhkp0y+sJFtPWPGvt4tf15Bo50FTQvx0KTgZapaNwQyLlf
oDF2sKI/4ZnVkOw5zyGa11g8B2gZzrohosKyh/4Ks5bYuJejdBp0+hq6asVOYAjkcgArGKt2ieSD
CT2OaMlmrRFnJWyCTsq/d5cjexjzYhwANSSDg2/QJTI300kHOWMbij4HxMZVixehBF6+YBRlLDxP
9B4/iIyQztiO9JT4vHMODvQgHhgR1NVqkFpIAp8iQPQFLjZpeuZ1u6NEj+l20Wy8U3EHLIbbhbL0
mPRcZuomZjn7FpRpXQckbvMTTgfLLeY0Mswocvfs8/uS2mIRYPEZgKoFj7syCFSdq/IbSYmyMjVq
F5/uaYrEKvrcojOimHSLK+yG6J1hVcNUMniUQkNqLEGGfGT656CEIHXvF99T5Vq+djSfL8DD86Jb
LMRJ4HFL1j9nzsDGcWVN68PGUM2kZfsw9sNG2spA2JW/Z9UujZhXw+RiRDzf0DP/40rsqfS/KYs+
2ebHxVyTklpDx9mInC/J61LPanSIEcnAZ+i+X2Ig32OssnBQ3DYJCp17LZa8kAV5+R28VZKNdN7B
ncI5VLlfDmvdsg14iaJvrbxr9u28x6SvgTxQVcjB2WVj+HnzG5yf4bJRFgYzUFbVA1AFHJYjS5wV
IiHjsQY7WWRCq97IaVU2vFYmgQY6hnFQyZWDnFw3GOEkdGavr6DIfdfg9+zX38jaKJ868sEFFQkI
vjIBtG7c2bEmrvvEgHDyyiRfV+LUSZ+DeM64vF+XF61o9I3tmugLCrZIlotHobQCdMadvKqb0gh9
0TsHvRzJZuVIiw8Dluagy1dDnDgJq5ceof7iapvAljN7aLvH+v7txNG0YV4DuIwEG5MjQb6qDJsL
/hR9SLNGKK+jw2q37B3weNQpV2tKrtP2O0GBbQbYdshzBRKVl9GFLXuR5N8D8m7CNsGx1w3F5kbf
f9uiDl7G2xdVukcY4GeOfgPFUafWOOFA6gu3VAJRwhqKtjRCfrODe+aoYSkTAnAU2BIueWVjCzDi
CP8hj2a2rfa6kr1NMckh76oyGzxM77EAL63on/+gQcthzlS51/gJ/9EaFX7Bu70v6towJKyImVNu
Iryfd+bwHqiN149EMWA1ATA0LucnQwLzda6DGgtS0VacDhzJF03arsZtCfEa8qGoqvbZaIVudSwA
ix7FttDfq3TYsplvQ2VqagyQggthTix9wCb6QMaGnWZssN50P1D564kR7P3ul7kWmp6mik4i7JMU
XlIMmlzd2TNVTx98QIgq7V5jgCDQhHJxAHu0fwBSESrUYI+6VLoZEO+X2uZrSksUyYCFPkN+CMfr
hplCPyDepDauK2wlHX4ky92C5S9Z39iJvfeqIcLcOBB0hwpHJO3SCIsKYqFawkU/lFO3DAEnsKND
ovsHzov+yRT7HOHXGPFnn3hsKEwd2bC98Qe4y0ebAUO43Y2dN/GQv0To3fLiv3LW4DgRe6qmVtq7
scl9RM2m2Vjx/3PuAwmHAFSW9FoG5Siu6FrDWci5yPODova0pcsgkBmSmWiKc4QrNf5FnlKTwB2U
kWqIzu/fMWb39bBB10tGDJ8aoRFPKNNWX+tzzUwVTg6BR5l0/GZRPwswUTGt0vkoQy8jSM6vKthG
eHJOJTjZ994eiNOVeXixb+LfqS0HETGk/eTwNBCMrkzM2tUb9b0Y8/BE5cpyrQSmjOtg0pVP65Ag
rP0gWA/zQM6xZZMDdjnbuvS7IXDKrmYuRgRZq6UBO5h5rWeTIudy2iQJJxka3Q+o6KMzbesfh9c1
1QmAHbIBv0nYGLaLHtkIXFb2chRKDw6eYSrxuDqbJfXB04/opRMhwLBx62y7+KddNbhDTZodgyty
zQmIlcDXEwNWnplnZ4ZZfNlaQx+n9aA7KDO0sDSDD86F5V4xZlPP4jT0MrMjRIWxoU20pMg4qI8B
IUEx7xOW3VdzDb1HuPsNrqF6VidT7fBqQAMf7idozhcxMalUM7KmW7y2o6d1MKqEbreaK+tkPGAM
qRtL9T1UaG1DtF0tdIbOJ6LpmB2Vyk/qb1Mi3Um4Go6UhX0xy3+OHOV3DBxAHuLN5u+fTpdB4htp
do4Wu08ujYaixRnYlYWaJ/AH5lz9wr7M8PTUFZ9rSU7ICx9xG0ynmrIGvfJWFBeHsqWoj4V/ulog
7d2t62xsE/jPyivqmZ9UjbouXyYGMYt+C2p6FVgNph5oTKjuS7UnkplZjkySEEeHxH6XP8NXSfFx
NE1y0/BHNtDQMoNpI7zvUwxxkKbaF1tWHM9c+lH67DtHoT55+lTLO9wkF0Lhssm8iB5HsiRHHl2l
DHtZ2PuYK4471v5Jf+TvaWIDsvl9ojyC/d3PycTTVWIx1P6QSOjUnEp4BDlG/80LL5O/BJ8YSsYc
gmfr0ZFO94RTCMZwocvdtEgNTGrG//5w3ATdE8yZYxKQpYx6pZ8+bqgmxo+DUtNpvAAR38vejNTb
XBbPLCKI9fuhmbGPxOjdmq6fAZUvMAhqFvghob0L+VkvPB7+FLiKHu3uceGXMY5UL2wGBCN+X7+5
iXqoTLSMhx21rc7WniDQqZeHBpHWypIYIhvFx3A43mlVHu7bLy/UBkM9yKTLGpQU75IgUlTse3QB
/BYle5h3ke/RJcP60jtRGDeCgkqAHn064mn05pwPT9vylCyNx13/FGtNN6MtqQSqyBoWK57fQ868
sbJx4J+0Lq1ndSRqYdca/1sAO746GTFmq7oVo+V60DZGoFYPR2Reau/uMbdwNC+8Z7ROMDOcur3N
fstG1f+oGhXOe92gbwyo6xXv6DJ/KMfM3MromOvO6XcZGfFbQTD8FVsPFMcyhgAEDvma9hXF7t8x
n2B03i8rmZ2pn4hk+iX/aYgQg1HpC/6CIp3YwrxdrsGOJ6cIFHHyki92w7WlnSed5nHfYcumeYSM
Z4rGCr1bNhBd0ryMfRd7D8z+NB157Kjh8LYNr/DZoAGRFfW08QTCyT73/e+yDvpH3phzu5Xz5bva
uFMyJ/Ah75YxwUb7Zs5DitfMuNq4nWQuQ+3vZjyqyaLVOFbGgH8Fc1RwlJ2XynULuuAoSZVYLObH
TQKz3IjzdGxkClLI3/AgwJaCfUJvFn2S5xip4AJQEksSG6D8rGuQ1ue8fyh11sRHqSyS8aB+zMuu
O+J1GRSJ/gVGy8/IN4dj5/tK3XquM3TsYZ5CwT+Oh12j/JlInUEW4pkiYyA/ieZPzmgavuQY5AB6
cvvBMNtH8Zxp/dskSBMIiES8gtuDA6rMmo0d2nVut9ZLZkM5zhilDuL6uTLE0bm+hM87lFNKVtn8
LtU7UCMCLPx26JXRhW02o8r8ANIq4p6r6hRWPbHtkLQ5isPwZcdFzrqHk6gUg/5RAiHFLrxvX2fS
gDdDo+QTwlf08ZZ7pPxyBD6/IZHvDGyb+goVn9rGe/IAlpnxPSUKQwvozYlnSSHDf0WQsVcgCAls
a6EWo2VKxdA+lkJdxF4Xf6wKWV2H1qnhOkSHRnOyjn/5H0UMs2JBUOgNh5tQYT/k9rssO6rWKZ09
SjyuXJdYNG72otEXQaqblSse2gRsd7+GTIFMwVu38+FBdYoaN8QJVcdcd1x2FsLQODuDxAGbGKD+
xAY7BfOeVhkO/j25EE9Ccvbk2O4e8uoKzAl867TF3wl5EGGy6RrUmn+frAhUkBOHkORC4Xh1ON1Y
mKNmdWd2tc7W0w0Yn979HBEFGlCYKJtn/NIzYQxGxyKiinCNKu+FG437S55qBwjyJCH0Jide4dS4
Mwdok5mDYyL8rvP3eP6xXCC6GhKcOo5VzcaIy+AOfaFc7LUEfA2XR6VBi7hbJNLb4W+AOsI6KpuL
AAkwgiBaNXl2AVU4VbJ3VZA5ar/9MMxWRxkVPhMnqferjXHCOOPz+VCryWel5M74jvE7P3GTuD3p
tFdYYqyNFiZD9vrew03tKFe8T8+z+zkArNgvEeayFVUfFjnj8zBqDxfRSb0goje+XLN6rbw3Dj58
IFNonSGai04vMWVUVKTu0wCrtFe6rYGfaTwHZloQZoCaPKOKsOh9NcIzIoR+5QViskjR/REZUyvW
77HZsdS3fuTN9qTnao2cXSex4eLYutllLmxPB8oJJ9i+ljNRTwObLGCrS1ooODJPb1KV7y/KnQS5
hKXLXnF/u12gQoCbbNx0Pp3zSQPKxvC0eYBQJRT4pMpSOGyrhZaZrrl8JHPm17d798bWPJnT6+Gv
m9WNY8yptEJrK3doJpvHrB8k6Qn/917PdfMsJ5hghKYuLsEzxxr/N/ZcgZTrPipGmDNvmei9cM7f
2pZIoyHdycG23Q/mZD7s9U5ribx93VHTsrUXyABmXFG5GOsjafiPk4DOc97+xl4t9XspRaj25uJH
Po/dq92L/tVHVKTquDSdxvvIdkAinQeFi1VwnVPgs84QgX1fSj2D37oFFzJi6FkbqNiA9n0mtHeT
Lg8IsKjhq6rR74C/+xCcQWLn06iHnPTJ7JMIing4i4anV2IWOZQNhUh5XZYiIi4RTyreIXcsKqpO
uHtG3iDm8YhExLNrpyl1dPAWBEQ2k+2TNBl+chlBwJHYhobTc8voSqY+hrn5ahnxROUncWiwc0oE
TpG510sBVAQbOIEou1Vk953rVK/uakCfTDXd3oKZLFt25IRT681MBf01WIxq5fb8YGZvfYopLuSu
hA9/u2eTthrl8wGIcWK1iD3kFaVeq3eRZJ5+6oH8N3xA3D/SM9vXdAvdLovjtTzmn4cjfDfMIa77
t+ngfUTzi6vUWZmI7laGtY+BASssK9qTuSEDv5dHPivJW/gjfTQ2ChcOjJ7g2NoN2Qci/NGcGU1v
fnrkjP3CNVbRkKPMEG4s6nJTCWrJgSlfmVkKqHWKgOkLSZCkm7NmrfC/CcpxPl+QKVD4rmXik1FN
n2lLjOjKnu2umDEFg0/cmStTjfFjgTKylG6MrjdnnBNSHo9CmQ2muz2WoeeTy6R/IGoKLGD+acNv
sjtdia3OfNCScKE6S5RE8zG8gaZ/o3ulMQo191qDRr9rWu+tKEddLCVdpFkX4CsEZ65uzysZ2fHW
kGc+KSOai/j9pupm5dcTebcj6moTw3CQucu/yeCXX2iGN/Ky8T6+EhempD4SX5dBGe1KhoGwZnKu
AuWd3ZRpwW40teqtYwkva4EALsHBW7rLfjHwf4MKZZwmqifMYcY3NIysy8/6aKn2BiDYogXPqb8m
ycZS3CLWZ1ELP9TdzMnBQG7vxnRzHy8BD9Ino2oIy9iPXWOfJQF7hYPIpqyWhdz20QkOo1eTI9hy
0S3y0a/xl5JhgiJFUCGGoNap8sQr2w9kFyVqBAaWWdDaFlaaes7z35KkHuWgGC8dW0dTr96u67lc
6F70yYHeAzIG3+8kugKQT2w7oic+4TpQ3dEPaPk8of2orImhnr38HVt64niYsUImfSl3B0v5SSnh
AkgMfgibOYsKvCmZpiVnTQx8r95w1P8QhM3mInBQ6uFQdSYUW6hkeFgc8zVrd+fj/wwHf5np0aiW
wATx2xUMqordLs/7qLxXugc7UulWgYN/m+kGouyojldlsZFTj1A0S5QdQ8WWjk2kejWrsyqFngk9
C6dHSCCGMflZZQo5GWu6j1MQmImPXtHPf77HrLeYl6T3xDldyY15YvJs1qwofaFjt7IDYEPl+vkF
HAv/3lBRJ/HOL5c7IsLiCqGSId9fRybHXOTd36Kx/lBQG4yZMne/3VSlJUcoRqqt0vyd/8TEeCE3
QN+RBb4+xSe7lXMqeuUIBGi6D4W1q2rqdw9QR3zVscn/JgasMSBbykD0NfM8ErpDmN5DbFI2CBzC
DO6tpZcSmc9xJKFBvvVn0KIiY7qXfqg2olHshbmS/3QIXuu5Fub/RxHHporKN6BDbV/pF7fd+J8n
r3z0SjPKXH84q0wkl/B49Bmok7S/1/VvPHVgR7GJTtpzVj265TdXL6WqFo0xE3NsWdN7nbzvJ+W6
oRNjsGsAwwTzaWM3iJ2oR1BbFD1MKImuVkWcxVNG9+6BG9+izn0D/QrWpeyvLqNRCyBGL113iCch
+HbkpOCWfl5g1J1uQlqqJGMZZuU6L9pt/iM4UJ5MUk8UjkYiZe/M75fXUlewvxYYNUJoW2LHpi/v
4tBqgpvZ5sBatn/iZAWkfI1iaVyJ0nVuIb0LVNUxK64SWK5v6bNRDZ0XA/CDiBPpGgyVVq+Yt4iF
UdR8qUPu3rIAllpB04CVaVTLbIkg7P4hTCJJ0iHRHFFaS459OxjQnvno6Fx0vw8pBo1H1jNn9Ed7
t5EMTGFloI10xObGkFlUuEU1jJJrJmZ6/gSFMOnD0Nwi7L738mWGuVB5EB+GGQYKKLg25rlV14kq
jxFJ1OyXwv654oFZfagzLJTyicJK8VgCeYPo+G1ogxrfivMb8ww5GWI/kP7764BvY+XgmWx/Ke0r
MtlYN2cmgMcV4fuiAzO3sprD4wj/AGt/XxJa4vb0ik66v23uoo0phOAC933Su2oh41LKikyreyXs
v5syxTEQaweUipwXmyzhvzQ2oQhWLwYsgoBhW2JqPFsEXWKD6EfIiwbPALtw/mpLw2TiJfGqrKSt
7AfZHMWy9BdLSvOnUejbyUy+o+OuRgVPIdqdd6v2ySAaI7rQ9PvelxnqVNlD+dyFr7KHkYq4N6mG
NZbzCbKgDpZ36G0Snm7RZ4AIF2OOJ1vWwN0IIurmy3Vdc+3xAfc6n7fkqnbj2t0uiqUv0fYbmjwf
lKvzNgH2R6NlFwQz/7dVeWQCu6GA0vZhoBT5DdfVefK4ZeyXA0nA3M0QwJVgGWs8c/kIWbYEkLu4
ovsoywmKvVxaB+iVhqTyvKT5n9jWc/A97HMA6WGNlumgwed6hVHN9FiT1RPUpMYpVmSqO1ZhKwqM
+HFY1WE7huYNB8PlHkZhxQsoZQuurObOzZsXybqppz0BI5YJN+TX8uGoqG5G60GiXeLPHtWi5RMX
BV58th2hXUUY0VCZYc/EHsxr4/h0ltDXU83pt1yMiS3ijzCqtXm92/lEzEKdnpDW0MUc0EX3UAs1
kxjhwslPPdkXZrW+7TRIdLFvBX1uSirlgCL6591qSTqKY145YAKCO3K6sCICFFZLf4c8QlcOrjo+
Cc+wBypxueCn5t4ZnneL/lZDtJnpEBapcepMzmqPZKpl8Rpp9kRlRucgplwamqMclEypEnZREFY5
D2VnQwHBc9tEv+S57YglY99MQNkRHGY62s1KiqJZk/01J4fgLn9EwkZSye5qjLtneFWSH3WRR6/M
RnNeGuHBou5PKvRuR4uEXcNEzJHPr/2/b7Pm+Xitoc7zZ3sFXo+KRQfnjmZBgmmZeJLba47IHq8V
zpabh+55U4AwcvPW2MGpkD5qo5ccV7jmCXFKFWCXRD30Z28mYzxiETU8nDFe9NLp3fCHbcHt+yB9
WLemmGgjawL99OAH/ILlCFbu/fgBS6wgFIPevGwoGhUltqop0fFXccID56MUetNdzw/B2oRVTwkr
stMichuDdfdXx/iA7cB3Id5nh8rwByKiRq+qzuZofb2reRjbfSI20WF+8iZN7FDM5Nw/8H+emVlG
5eodNxmwFJrV9dwH7deHyrGCdrWal+efI0OkPYca0fSGyuNgCeKWlJpAcXzfl7DlkV+tr6u3Apbd
lpzHlBk1dpqMQNsHi/Z7RX1qejvoNI8sBMnnH/wnZSK2K67LTCuFHUh9caiyFVIOSXI+i0VBUJ3i
wylUcr75BwAHwS1LqOPMBGEjzEF3G0d6Q4EAum20b6M0A+x0NIeoR/N7RngZl/BSwzfUI3Ts+ttu
ViAKBmTVQIgVMVSFxCatK89m/Zshzffl34AmLJnI/mgLtRl2jNzUJMoAGZpa5HakfCd0VfuztKAi
tZVTj6E5iKTmGEibMf/HhrtBmjk4uUsjniSRgAfWgTWBT0iVYpz482mUf1X32K1vnDyIFM8d4kSX
k5cGrGNJXA5wJzaIJo0R/rggfcr/6xE70HSQ9oUZBJwqS0LT0V38nnIYQxlIMKvbTXDBwpN1kDf8
/XHA9E41q7dbIxt3wPWQQuFitjmu1GADs/EHj/gMzSn4bY15VmCt/cZgUqr1CpjUh3YBDNhSeb2Q
RknfWm1csctNHiy5QbVwbWQyC968Qh4JvNihHofbFc/lkZTsaZeA++5k0HNlNgXQ1KR7qO/T9bIM
9u9Xe800BuKgI7EicGGy40TFZZ9VkSE7psuQw+9mVJhTF7akRK+lYDRLt1GTyPV+cKHZh3VVALkC
RrHgoDBc7AO/MZPqnjDpbwOyOkOea6LWPgG6bS/wtf5VjwWt8hsOzpxzuckjPeN9MhJ10flUpT3U
CjAtkDlIO5lUhLnf5ihUjGkT3bGPo1NraasuLJxQFhaY9H6pxqCWSR/as44IDBqVkmo6e4C6GCRt
Quhts4oZBECCWtJtIDp5kKsMafJ58OIIWNvxUTu5H1/NuHRBZAL6U3No8aZiuHIEe6bius3ocZA7
IajMQM5Bh7zd/OIo0kY0mAliooDWhTqDIq8AmIrGyax1ajZp7sggs6rS9tJRGNnDPCUoEsJC6coZ
1rtrSEM9yTrU+JKzLXyPeFL6zjyQWl7qTpz9AL0ox47VeXZYgxsRXgmyJ2ge20zc4tib3nvbkkLG
qU/MZnhdvmmRGdAygLr7++eMFWMtyvV680dGG1HCDafgUvZPSgyLwjIE7NjGWNNF9kPVhNUiAPyg
g+JZtdnEZ5mFCsYV+0PWhhW/r4aBksud5WszDfq0WKEZNqA7KyhWhtqOdse4qYzapGslLzi0F10G
W47HYAkxUEHwBmczWHqjJdpbDobIhMwbHRM2c0J6vgOoETJhkPrhQ+tSFPUDKXz+QcwZ5hQ3OOY/
fk2hItaOSZ1gNgmPtD4EL4a/tZszxQQYHcuWOD8nVF2Y0u1EmuWoVd5e6itfz7W30f/Jy/p4BDiZ
akxvgc8QwJMTbsB93RHvmGBJZoeLkXjVd6hCgQyqgG1OYRdtVCghlMQ1oS7XsdO4IvcUJ1jS69jM
5Vs4O9Vt4T7FFoj0EzLGTOiOscMsABBopleVvq76Y0FOPi1AY/+a2K5znCpwdsmGFlNIGOS6E9Ao
ijxhniTCrd/3mW1/VSyHb0KSpgapkhpDrgRBehuIHrGxGBkXFwXE1RrUAJkp/BFzqkM6UVMww312
ZkEUf0RZqUBkniV83AgVbDP4S/wWrBOs8NQAzdf9glOTnv9Sy/Lf2v705kkUkCClMbLeFHzfwL3H
933Oe1zqW1eutSqD57m4RQ6YjU3lbqVZ6wi1PpcwOH4n8GNLwAY5n2LGQprThDgw4bYT0Gi24VYD
j21iODAcVbUqnEwit1ltsFI0azCsYPT5r84zLCF+iHUr+xqtt54D2EGd4u2LKvLuNzWJWrOIIfzm
4sjmexGkqrBGviVS1CCRB8bYqhknhjcErwPuHK2C6hfTzsaGFqbtR/RQhXQnyRXv5wgdfBSbxD3k
/4b+q/qtIOJC+2W21DifFzHud/uXZDXqvT4SHZ1G/IOWKetGM1XGdWVmMC+T3+vIvB72pmQRylgY
Lm5WOSWDme2qQLyFrky3HO/u/Jo862swfMweHSK7D3qyC7xsWRPGDX/YwdkqIl7VCSS8bvuHNDkG
cFHclpaLkbfamFBuIEcocuZeZZrkWZb+TEOyxvwjxv/yUOXv4U7XilIiv4tusruFwpUI/lD9i/+z
P16JhLjsEOwFcXk/Jo7TQGaCgIwQNmfPjgPWB06TWL5EEh4pDIVgjMUvJKdvu7aYDnWhptg+kBFa
1LtKXTNGWJBUrt9SEbbigz1I/Ewzo4L5SnhtAllhRtAwVQ0F37Atj1vtAEjnDxJOuLvn4nNqX2Cb
wmo9ujNW9zqokaOG3vYDbUiybLg26KbThnpaefE33394rkFYahf1WBRM38RTc8ZaK/X3tyz0mZFp
yGwHibkM9BoWl9nVu4T7qMY+mY47upWeZcbf7d5Ex0xNoyQL+jlH0f+3oYTliogOrWVSsHQwc2rQ
VGzHgYsLMpRhKxPAjUO8aHvIwR97OluDGWst5FhFeD26gjCZ/Q/1bVHIw05+Ug1QxAiW/TJukq7y
OkP/Evq9rSGiRpsPY5+2BV5TNfvknY/izQnPmZRI881dlu/XQnlB7+q/vI4UD+oGfLuUw4bvNdKQ
NisVTr+XuQQuvqwzvkhJYoNYhBufVdfHkrl9X5iZhfXaFZ7THDRlHk3lpr3bLdZtyNyTmz8+2sVO
wokgh/R6wx7EjQl8W8cCKUMSveSLiJ7iZkTm7Qqp9AK96FNwo/4kHH2tphL41IwHmBPBH4MmrqHU
PxJKzl+pu7hVIe1/T9UCNnxgAnBlvQHsD9pBLP+xlGv/hEyvrFsJE8fBUNLGSUDcXiJTjMDq35CL
XYMgtqy6GIVHiMko6rdD1ROrpyDnVQctKS9xC02fJ1RNNowWn/cGkEX/Pdfd7FEJeKeCiB2LAFrh
agwYJXakXM4fW5USgaWzCt2Yty89d0y8s4D9VJIqJ68vdQaiYFik+EuTcPjjfyBkqtQR8Fmyq+fc
aD2375bmoAyHGZpz/qVvFeFVQmWi08QGtYr+Nl+VZL8DzBAuR/ryx+WR5UZa1l/xc+64wrn6alRG
sDJe8mJYqfwq6dvix7sCAM9xOuhd1h4mZOXRfFu6HREqvqZS043IAiTtFmBRdmjHwHpO/ZaVWett
PTL4wATHNy6tosr3Loejd7c5Ktp1e3U1QUDXDEv7H/SWzqPTL8bD7sRDYalq5NEav39y2daZE2S/
CNaygVhnZ5zvIGlbcE5y/2GFRTKQEkYokJXc2txSQ0w8oyQXM4Qey//0Agkiwd4K8gPEmBqcek/g
lqVo/qT7uTk17I40e/y9BOZ6oCRQtysGoJ3jPd/OUV1rO+QMoTUvUHnwPau7CArHEyYutQe684aK
Du82DrkVhQ+4+lE+TWMqdz0NYZJp+PjGSd7neYX639Qb5CP1BJ5AFUbk8aHYEuTmilIxlpXAD814
mgfZN2xbofQ2+x5sGB8iiHpXU8p66icfDRoVC1wIr8aYjN1ZEtcZ17gXi9TYLkIhqFZqjNX6Su/a
DRSx6UOSNNdfUxVLgibGObie6qeE6VO+vgSobdajoLebWHGJ8aqc7aimbtjaI98HqZK1rk4yB6Dr
8cuo6GZpg68XePW43gmRxro7mjFxPzPILZs9XDWYGoSWFpCnS/3+JOZ2+GUwMgExg11agaUBlALs
TBd4knSRIlaK3W5umpjUE/XO8AuokXkO0H2htl2H3fiY+pgnHA61eZb7POlnKE2DtoLrIP/uZYV7
OPFYLhVDQJZ4zt2X+74kO+6LE1Pwoizur6cRN62viPlQoq4HcQADawYsZbyxXTIQvVZGrbFZp6o7
WfQiLCqV0BABCEDP77OM1Y6hkCKpU5TDHmxOHYWHBhVlClPowGB9fB31s8wYJ25FVz47QdzRLS/x
TAi6khYLcCGey0CFOEecQAg7LjmLtcZQoP9RpD24Sr00ZXmptmWOBQo1/5rnyGeitXaohQJb/NNI
ZA3e5gSXQV1ILrNim83PCmyqLBQ1gqKrtYiZayzFaYN0gVnNmHkt3Bu+xOWb1ji2X4LLnc20t7Ex
aqq5jW6YI+bWxJdT+W1H/5J4+SoAL6FeMW9BBnA3UQz1mjuOODgT/RHECjLPU7H04ysB0wZPUkkW
7Yq3LyENXIqXqLQ+UU+h/kiLNZelNu6kvT4DBKsBtkKmoJ+5n+5G1Tn+Pb9csskPeZyR5DEeaPf/
tzyZFx9+HssyECGlCFnFFpg0irQWFxnu7ChSk/6fEDSU+48sFizwktPoW0GiesQTHJ/LZzFVmC+D
yVypuNEcxZ1p9Kyrvnpva3SO1dmLYyPCXICpoPdHS3isH1S28BqRlK506RZkctTpyBGpx2mITL6D
61F8A2Hb+YQQquFoDAeJ82xTsn737WnKWYQS8peOyRC9MQKiXijc+OhWt7vyGqY6uNgDSeSPeXrs
+C18ZCKzk7Y8BHykp8gv2fal+ZL0LTe6DFy5IR4KEhOD8o1vIeg3yU4sPTePAw935GU/OTZlnUHG
j1onX6wpToQdXKaOiQWiN9d0Yy4szHhme0V5vK0+l3vtT2zmm8OQXvNvgZBEFq6/zkYPF/OWruik
7Rs7+03mls3jLZxi4nCa821pP0aNoZABNzxoG/LD6qvXx3p5PPC1e8g/Xapo1at+RlgbxqHQHG/B
uaeHVzxQBsXgnLw0x0jvC8RK27vrw8ooqonn5p8cGTr66vQanJMTZmHxqz/uzYqN45fnFpwuZgGA
p807mlSgdggzRy5UNNrqFu27O3tn7Dw+Z7BzPGgli+0yM/j1YOJGUFW8gYd8o4X6l8qNM0j3hT+m
gL+9toS2PF+P0suUuBHrsmaHP/4mAQV1cTNWuGpkela90GlRvYZpfFd4g96sc1EZeqk0OvDbaVUG
Q2zSBJCjVEksuk+r8fEl+vCV69d9ryJCW/nUAEKwwhzqsYwfbHvT8fesBCt9ycCtN+YnpK/8reY7
1c7BvX50j+/UA/7SvokUtOqdHGVPzXIYN4FYk5AHZxCjXJJxEf6SYaLMiyOrKvwwX1BaGxcb04/z
/hPnbD9/Dk7UJ/WlBRu2zW/RVU0UwGzhzLuH7NNter9cM8/bX+A/adr/GWdh4P9Kg3IQpvCh60jm
hFKMzMOkxLUFJE/xnXG/ie6P/ybYUn7/8EQhkCyEjtomHHCxwcAGOdvofiAUDLGExJsMzNU2MDLY
b4SQCxFDjJSrY7tzZ3yUNMjP4niOpx2rqMbK77KwRvKjb+OcbGtabyinQvBdGuarPzUT4+6MUaiy
qInNZ8KCHMdxrGbvv5a3tvxiS6Kf9x/UhhNlV75rzhzwhd8VKH+feRYwPTF1WdgX54KPVflMG2Oi
waF5udN/AD+l4pcsR9a7khMEOR+N45koy0YHBn2o8ndy8AWA7hnNigqDJfwadBWyprVhaeNlPme0
0HWysOJRIoCvkazuoAbiTsBUQ3oOnGZ62GiA60S6UaMRIerhj+4S2AOnFXDlzw3OYoVP1q2S8lvA
zDiNvRtk8XEOQ2liYbbT8T7gxMZe/gFefEtPWLttBxBduSgrz92t08aTQENHRtPOOPhQ6Ey935Xi
YLOd35gPG8IxJozhMoXvKwtfKaaqD6iRsjqBhvk+BjrQFhk+E5n2VIO0f5ufmMG9l+dZq9aJxdpE
PVP1GVD4AeIk/mHSQ0imoYwYHcOqXYb51p3mpTDWBIaot5pww08HeEtRgAJ+E9VhgQrNZBb5BB2a
gCxc7oOdmb2Twj1ea7FMVuoB5yeplp1q/lK+rBU6Pez5AilEckEdojzvnyK7oMFp7ODnvnXv+PGK
bCQTDp49AwT2rGTn7TCmVWPfpqshQrtHLH5+zUkLT/AutE1JghAOHL92S+WlIP/mUKH2ivsySlFV
geqVWteeNPXg/z5auBCtCaBT/QdXVAKOUXcY8ORZLaScdH8uBBVnrGc3txqoq/2Nz2l3fa2f9vyf
ZIbvUe75kxuwgVJd9smyS2WEF765Q6UpRM6e2d9g2JYxTFm4SMXWDqs2FcKJCTAM8+T34GPq0Z/e
xG7uIl89korz4hS6JBYtkXLNnBGOwwOQrAQdfH2kOm3z25KbmZWVURNYpJFhmWVcpatl6OZWC3CC
5xugnYouEoZuCG0DeDsvBvU8+vvj3d+e5P0eghEuE00EaAx08ahLTR46RGkUAMRafYHhxqmmEVTz
udHq9IgUCsS9ezxBV5BUZVxP09qRVd1vjkiFGj1xd3rQY9sWIc0AIkycLgN0/mB624JNCO2soSKH
4PzMIdi5V0kx7qzHADHltN91PaX+7EBo4BH+pmb8EH8N2pdAr7nzEZDDx7DWPUM/pvGWgCb7G448
DELp6c4T41Qit391tW/DS4LR1P4KbPd0516sul0KxHm4Rn3ABeCMkonycSKNGLc94OUYYpKL9Aui
7Wk7umD6XFkKfso5nnybWFz/D5N9Qq5xe+CP+m18l8MEoTMHld5WxdD/jMOb7gStMCOJG9IvvtqU
p4pd64pxlgVbs6whPbBC39YOPLTEDZEinTCb7gnUKDiFh29QX4sxOIBOyop4nBeohG3uuTzBvSOE
B6dnRFsgEX7pkL/gGkLWN1nWarLRhr/ChzuRXvK+4XAd/8hAtnJFKea1/r6coRf3s+Xq/j1pQEQB
muLhTrDVFuGeoO4f+ksaqbvOo6Oj7x1gA8hCom+QWLIZtiXRvOvOCet7dPAMyWfarY0M6aVT0EIM
GGtpItm8bdFDAw5XpdTJpbV6MNUbCxbR5QdI0GzAOyh0JzNG/5G8vGIOPOXI56vEKdi8HT3Y7h5G
iIoRyu4GTImdjS9wNYltMxKlxtcdXQdzOJfRsm45mXMBcnbpOAfqg6U6UzZWb/ioW/C5rg7VBIHh
4Blg9vYLue15B41Shhb96Zx0zW0i84Es8VWmUpJH1P9o98fTSlfDzFNONEJ9nRi8HtTI/WkDDQVh
+c5Am2lJ2G95c980o29FX0tsM3M3kfKTH/YFxbjTlba7Dn5uw7ulio7bc6IMj8u2aUbNFYl9H6wz
eMyXFl8wKhjIxzav9jJ0m74hD5y7vSjaC0lI5Zcdj51m5XFPWu+zl0M8An65RH81OYsWQX36jXIJ
ARBKBjTP2h5hVU2hY8ZBPd6+QEBnvCqTZS24kqLYGYketi89GSR/INEGhUbN5soMTF0BSwv8K/OV
pAlerGY3o3QNl7RhJN9EmV4eg2Zd+fLFm14k4MibuM88FOoJinyeowcyt87qKiMuLJMY77hMOxoD
/23QRrbco3NhV3BpEYrfgirXZBeofNh6j+/sDEJ+hzwgtC/KjU/i5c3dS5A3/2TxGv9mL8K6Y/is
ttUUvqVH/mgoH4uHfJ1HRhpG9drhPe5/ZJG3LUjC8Jcgn3Bv28/NeU3G4+yszHVH4ORx6Eb2C0aP
oDrLEwsHqY0j6q/EJ8qOAxR3QZ0VK9dTWXqICa2QLADfsnD5BGRbAuLajfwpMlYfOPNuZsl3Bsdo
l8iUKTZB4u9O9ljrCLrk9m+aUazMG6BqcO0Z6JEjdQ5iZnP5FDvUHFAg43XN/bXU9HF64Lt7KXQk
25eHZ7/lcaTPwPEkP2OXMxOABStd8kQcWBzgsVGEzQgZMC2d03bMpSTV23FX6cDjcHMLn2GuMRSW
GOXtUw5e2PMw+o32pN4L2NwhJeaMdRpB59136OtPugcttDlW7IjZXxjjV/Z7ea4deyPFeFk4bbmF
B4WtXVcTOjzrZZyiST3GP235luRTkKoZu/Fdec5G+nbjA02c4lgRyAPesIEvzEJXc8BHGj7m/qvZ
WoXaubsWBBSlHIT+r0WvkvFAdJNKnQdg5rQWlK+u05f8kEXK03H+Vg+gh91+S7KzBsOAgQZlDvKz
R3CjGI8WJjAuaz6yrtfIwZkDq9vJOKO2xqif6MuR5r6+BEc8pXxj8MIWnsj53kiqTcJVKBctJKqn
bCHQzfJ8+IeIomBxS4y0Ohodbs3qZG6WnGQ7BlUN2yI7ZdeMYnfne4nnkN8xzrvlNqwm0RJTrCDn
iNomjv9h3duT1Ia4uonIZ5K3niW5qED2ABwJUjyaoAM9rqJGz7DrF9INlIfp85olGjx8OqeXGYD0
denAgbbrboOwFF75jBaXiubLRSuyeK02BdXnQJpIwszXRgqqbKzGZpQqujxusuoo47wMrfDy8ayW
cZTHL4TxasI3gnawaFQY6ooeYFTp8i741CJRiLOQlQ0f0HRR61RVq6bf1toTkhgH4Gp87hU6Jk6H
3xRvZ8KJ2Dgxeolgq7iTu+8/YSwYgA/BVePfm2XhjKuxtjN7mzhDcVf9JFnW8wRvh7WsrjS81Y/3
jqyXqxi0dcCniQ+9txpXXlOSwEw4cQK5hE9i5ILMntYe6O1bwJITL9mSIFaylMFju8Yo6UFQgyZJ
GwlvwJihUo6mYeNTzrXRh5h1kdI6TjNUA1dR5XAaX8OwteIN8pvYodxR7aJGrsTY1z6KrFnaUlhE
EM2dVjKGe/VMLOzS9a7JVkFQAnvtzUEHSTPQ632ZiUqYttGqiCkPy8Yjrw3pNw7YwhwO5dE24Eik
Al7YgYB5sz+X3pOsjNl+v34VSQXh9iOa9b1AjkhTYd1BnvTDFmf8rmxTveVLSmg/Kb7INIBtKT3K
yvz94JgTBcXfeYA9vNb2UuBG2a5SanrM72n7/rde1EnIfTBmNGebTe5vGT/yyAefou0TaPLpQFwV
bFqD2qnZPSochIYEfEf2Qzw2rdIruA0SDFrfO8e5Lo1vUrwN8IkvS2MUgC+ZNSyHi3EUVigYAgf2
pNgF8GmTL7gTrE6JH5PgGmjc3Oyzuj3st1BVyYIxQ46QLgclMgMKyxhehI+pDcTQBqAjyEBY+/yL
doORjXlhD1Y20IOpXgmXkeK0Iz9E9Lu6ud/Ck/IZgjZyPelbLlcA3DN6r2tqktzEzHeZjZ6t6Z7k
dBz7Gm0m8En49Zg/HRuktCRBHiBI9GXKJmXWkOX0mHYK5dYX53dxIT944fVqrEbxhW63sDX1ygpb
Fni3GsPtIINbkcOByjpdOfT1jMrErNsFHVEt8rZH2ah8D+wRYFHjRBRCxZPg510yhy++5oYiYTkM
+4wf4JRxGevt81tycKBD+4QglVq5V31+iYr+8yJnbb56gmNVv8KPprs7PwzZ+7rl9xSb2rsPw2J9
kuy2jLE8cW5Mum9aSSU+0F8MK1EUzu3uxy3huEqwCNV578aU/HgKeCDIOWu7Mm5wkx6warH0jRkD
R6eO3r4R+NbkaRK5MIyTTJwh7+1yYd55nBtKWY8Q9lqCEEaKJ+iggq2SIJi7vmXAK7EANXw+5JGI
hU3xyHR5W1WggbpVnB+RnHnthXEA3/MHqUMYv249lJ1ksSpm2QMYDGq8lOGICYB9yMoM87SLZP5j
tOub67E3BiLi6NJR4TnfJjwyT3LBJCavlqxrE+gQdI5ggGjsW3f0qyTFpstn+taYwidwPFsJAiBH
T6egE9QT+v5DvR1Fwu8hl2vtpErjlczi1rK04/DM2EDY+JO5BoiVvTOYZJ0JhReJ7JKeDTnQa0JA
ebduu4qXtHcXC7MKatTzhh4i/0pY5LBxRiF1R6/fCehcDXWEizXnAMYtqfO2yHcPGdcioPagfB1i
9++8ncpYCB7spHlOII6wKU3nYoYD+RgfMo6y0gMatINQ5Smjf31lECmRwJ4teixJNpbOp5hK1Qmv
r4N5jD+5i6lnJqMugZP5z6rOKJ5ErSW4DWwd6Zg7BF2PoHYerHT43p/LzYSksJC1t3J7TBYDB2k2
en9HG8AC8rOI+TUCazbX+FoQSzxvnphGPvcTToN/Rh5yYgBXCOONu9W6vRo2z0YscFCIdu+tQ5m9
QPVHsy/Iq9ksy0V9uoLY+AmEaun8byeB64+Q+Y0IrkWVoOI47/u6DXxmFuW2j3/IayWhowai05tj
ou7fuWNwUZpTT1YEM20rP6r12RojoPeYjRN98pEQfMgjOneSk8D2u7ofkn6z/uayE5sR9fIzER2Y
8hMnZ/ht0PPGQzDfrEwUtSt8fwxqTGX8wQhxAMruqAnVmC8yItBtY50M9f/pdfDwNR5mihhvWhxI
9xQK73nJ+jfTr/CmKk2GoIRYywe09qlw+ZlXxMgYGZRz6Jx6HaEzNL7wS4MxtG05ofr/8uYAu8JQ
x048iRmA9RYtpKfOTm74Ekck2ZskqyuisMZOvK5Vf1dQOanjuIVgRsFVT5TBGbFnljSQ7fMdA2mx
Ct+NxpPR0ki6SbDXt/VoQfppMI53/LZflGK8HxxlFhFKx3Zk4JJWcVOCILqwFb71mDTnGrK8k5KK
61rR++OuSpRS5m6eMeqB4WIwjrYDpV6xYPPle9LEn99WMcKoqdppSqFZhEVMlYvYy4mXyasoAzjd
WfhEz0+9nFhHcHBg8AYw7VXHmd7h7dkONat0X5BTZz5oKtqiuqvXaRMcMfwGwjqnxhld8UJNHBkK
fYnF5NZ5cOxNpCdWFXUQ82yu0UVRgJhIdZsG9bDI0VUa9iSFr+XafwSaxmhsKou8d25pNLqp+7FO
nZjcnvPXLecoGMYl13lYg6m8WdmZFi+fusv3NnG05daSlptIot7wDw7L14YPRi9SP0LjY1Pz9eWr
JPUZ1HeFv+CLldjWMFyCOZGKdEsZ5QQlVZN9NjY0gDRRJJ2Jc75yZHLiqn0HpM+Ph5jJ3tHblpn4
y5n/sEzRHl2KWUGKlUGMVs305UHYoypBOJr3U+JJSZjdLqp4mVCrCjSXDyHPsrk3BBeEjxAYcy3/
Hper9ZfAftrbjaCLBHwzhIOyFPfELyRHlttraFNK0xWZF5+Jco6ObIdZYY0pqgtKXOwA5P52rZ5f
yJrxh9BD54+I4ARxulC8ZfIiUUhkEs+xYuf6NEA4IMxUNmaT0u/4+YqcBoU2e3BdML9TQXHF28Mm
VLpzy27u57LaSJc8g4gUf6kI2mwgwFDMPvOrmiqxV6rlkcKJ0T5KiAkEsMNdwZ+v6ZsXyrLRzuL8
W+KM5cjPvrHS/WF8Il04aEOhGPkhq+HDKOurZ2R4lvYnTlJlbIxzmdxKeheDMsEOzsSaTa5skOHW
lTr2etnqySY29LIKkoAl0z4zRpvB79rwhUJ5MHWCVy2F19TTxF1Zt0KD4aK/E4BGevEORyrR8mYa
6UPogxN8Sp42Th8cARagAQp7YYcIg61KI6IXS5l+cFuH/uibKyNXenh2t/0JBfIn7HuU4inxGwEg
RwozV/lr73P93Hl3hbnQBus57Iy+9dbZHw9HCYsTTMkgiALXK5tiJnSf1+fELca8c0Vd45CL+lSr
pEjJXqyYNtkb8mSM9Myhb8fXv6zI8iaS+hQmnMDJ9/HPiO7/CRepMBxET7nTYXy32mjoDkNIuATr
JmHZaRc6Xx4ozjQrldJPS0uHybyLGa10AAspTT+VY+NxfaDlHLDRreG5j39y7Tsg54EsqlHmNQNQ
XaYgAD8iCoQfTNy/Ntqn3gXCI8rJf5U+RkW/tbzvMTDF4IsDzAw2zQ+zFVAjgBd315U+XV1Nzus8
BDTVD/9bUycr4TxJ73H6JNAOFr9j4WaJnqUOR42gTVif9bO8M/6JnESpbqHuvZiMQvynC1Mptgio
OBhUkMpGUkBc2NwmYmiW7J+dyEx2g3oW3cuMjXhfTq+Jnk2QfjcxvqtK/vdg3pPyQ+7sX73AjAzJ
gBGCgPN/T+1eVKWbn+woB5cjWognpCMpdqJX1YI9gK7QMyccXeBCDOetP0/d+hRAUx+qgNHPZGBe
eaqsk81hUn+sumymM/45si8e7hetOBqyHnIXKrBhyRTYjzSrBdQJl8273rHW9x5aONvli0q7f09t
TF77i6sMBzRNkEwLjbmYZmzb/mn1U4mpFz/FuQCUUqA9zQGe0U6nWvbxLyU4LSvbmjYuM/vSbyUg
26EIh+uexxE5jjGqUGpsZ012s8MYohPGP6dMCTQA7Sv6LzQg7X8X94kZLqjiX7OSfFlUNwMfz/ir
0QWR4G3of6whgG+e/RsRGtyNP5kj8ij8Q3o0wrBT9Z2jZh7LrsMAR3R7GfKaEECY4KpI+DbDfIOw
QyR9rQ3Ll1zbglt4sD0BFCG36wC8lxeFFyLWi+mzh5wsTxdMkDrtug1QLpAYdGsYEvVXq9d8ExQy
/Gpjhda2/AR1MFzbH/9dn/3tk+jhbtuWyWhEk/5TxJLdkek0Ti826WpIIMemLmqBDw3FDQGaDMTE
dLEOFV1VSJgnjk+rmqHoCVhjW4utqbGSUWHBmH8S+qmCYuvVvEqX8LCec5uMIOzOiuzYNoGqO93e
e2EJ4j11XVdjTz6NcH+2eoZo/9LogBAa5VyyWoqYBSdC7EYmRy+dZNC/m+BgdgHYpZuQZK0jTVZW
3EntkbDxiur5R11Fe7jRP5r4yPIoSV7FSjCUCu/ekXV5Ky5HdU16lz+xwk9zwExvFAdZVClTZB1+
kAAAYodZIarJ1OkvhqVHZ/BjwKwQQhmQyN//KApm/tT9jMjAT0JF2sCKaUwYKqd85wj0mJPza0IY
p0sgSN3oj3SNNO7RMjjpCUhX4MuAt6TXKyh5PU8sdBgzU/2KEp1H0EjRnfMd8Cy88B1AK6gtCD4M
sTjkhSFsQhl8fl3NdE3Av1PAo3h+1bBD2OKbcwMi+6p/xKZlQ0eNm9300V3D4ZUvO6c11Wu8yfSy
BkuWI2QTBAK/S8Zy2oMyKYyXogy2nNzYY3O0Nhhg16ZdJ9nyOj6TFxNiq97XXQJxUYHwVveVi/jz
CeYM74DHII5TkXT3APLwRB0bUqtPIlNgdNin0MOmO7CGqbeDn4vL4Q4mLSJlpxIH0Lb1lVVSG405
Z2CU3uOp2dkmqa+l7QwK2g6C8/o2ueIFljJJKY7ppbXhAR21sm5m58+g/558BZaeiwnr808HPqTj
WmBgtRe5gMjoVtfJlUk9khktvXrA1FI/y4CHPofzaXqpswEc0nZSFsaH1muFps+3QtB322aupYHp
MMjrMsbpuOGOSGsfWuGzF5MY4Pm4/vIEtV1Sx7kXW9iS9y6yfQ384eFq7ohN4PwRzf56lKU6IK4T
l3nZccZgfp0TujOr8LK0P8RjJocokIHSgV0dDPcoq3bWfMsOHmxhnyiyIjcHof3iwNwVTV5W5jCu
0mwSAhKkmUFAiLh+KgELWSvbIaPai5aXAYL3wnqhYeLyT3DcOQOEWFW3T+9kxXkOXp6j2+Yot2jZ
6ARmjrLDBdsdlJ/yeeddbMFJom+6UmRzN3XsGCLDTMPcdFvX2MoujOThp26MwAX10m8xQ33tGJJX
x/2Kq/wp4C/K9t+UlizRorC2760MzzrMkRnVecJaBsjXZF6v84vl8Rsk3MYFrDQJWT1btFauYNbz
E8DhemVp4Spe2nCbqcaJH8KK38y2YT9WPPcgxP+6tSEEaTJ05AFUoA8QcOuC/Dhke9wunBnmdJSq
R5GR9gs+COSYO8+5QGu2KOkc7T81YEQoemQQXzIgiWqg07MxZYoVDkTKRrruECGkA7WqPk2DM45L
/5QxEP3od1rktaGmKH/zFeXHjF9/IZO/LP0IWkWny7H2hSPpPLUHHufnMdXlMHKyHaFQ8Xg+L010
0EtYCN2/9lgSPnbBPVVvSdX/hTSGHXdwmv+l6qV+vmcwcpb7JFzIDG2ZtAZdVSoLrB8UW3zls6wJ
Adyh0lqe78exbrPzxpKuzuOmCj4nbL02Viz8UKw6PBjUdNMpTDSgvqD74x0UhSGp6zkGOwDDeTf9
OoR+g5l2Nl3p1gQIHMt3eWSmQeveBozxHugxa8srOv5OeUnFffuBaZn16JFUCgRX3IO0v/MCwRS1
MkTjofBV+EYwzk6DNKu4Cx3sd+rSJsr/DBBzttKPn1xOoCYDHo+U3auLMpULw5AXUPXwXUtMo6l9
C7Vuz/I2hKd5xETtf2/52BGaEAbIdJwg8iHQkyR3aCcNU5MrN3UGCwoSwLjqEJIJ67bX4XSZwSWj
4HgBSOM5gku5E6t3HPJSBBNo8Cwg44Dp41uDmgzgI1NeHrfHjJhKvfKlLjqJgM+hj9J9Y/iDt80g
+hCcMxXaa4fTTRCXQ2tnavNlp3nqYAtNCbYtoRWetaUl2S3Z124SqkR1sNlkvXpc32poR11kxVse
itAeH+9/0J+l6I0cCKPLvFgrPZqGVoRQmaXdr4Yrl4uOo+6y8oZJZ+Fq+mN8DvnoA68VEWN+6QC4
HZv6gHBwr63SdMgScdAHQxzqts7ekBJWEp77iQJzd+D0Ex10aDLtqsYBnl1HeyyIrV4vXG98bcJj
EOTQh5vpyDxJE2PgqOKQ2j/i7M1faZGE77eBXgzmhwXjiObbQuRYkpOz7p++HXkuV1w/jX/Hff5b
LXcAzP6KjDPKPtdnob2SicaGLB3cB7nkmA2nX8kfEx9/IbPK5KT2dcu+gFrDnfJ590Q0s+DzRucJ
zrdgx/qFsXws2pIcVVvIlk4NsLzCt8yTcIz+u+wv2F/PiGJ3ShYXP9PTXTtKmrZgr1NSFSw0y0Gh
aoj9DsAfW8htfRsksDMQHA6XFgqIxpLUpKHKpwtN5MMy0o6O/c7slLgpzbu007MjpQFV/ft8k5F5
pO4c2df9mTvDlvQvzU7d+Pfgcncx21hLuabQWWYZ4+DYlRcYWNF88kXQEeZmwzoolxdgoL7wMrCV
UpcGlxoHl+0wIvnRmXg5Bj6A42VT7F6HgWgiDohbmWwV+lBv8DKZ6FELVXw4vYE4JM8nNThbcSFe
2yh9hvN6buy/oumbE0gz2JQ/0W1+dn3bEGzn/wJ6+v6O0Xb20fAXEd2bO7CBFIJ+pa9rdTKCZ1rI
ugjWwon7pM9+CzYUKYob7pVgxj7z8AOgMQ/rhFbie5G9Pv3TFR88D2scsrnlpvqx7D5Q73fl3pmU
5xz+n/f1wO4m84qlOsO7xvLgQWrOVHNGjlhvLqYF3+ImCqP+voGGOoqz7KPsuEanznwJzd8BpIH0
ybrF5AD9GlrZK5sJLwfgrQ1FLNweb3zywdiVVUljVsPEdhyYnKY4b3FGFOsjIh2zbMMCbhQQD4Hf
Hf+dJX1pS98ujm4jWDjIntsKP0kGED6T1zzVP3ix+MKVOj83WZgdMivoH5Unhcj8vKIQ7VUxciUq
xJXI7ZWAj31pghvBnnNg3TkD5fxshwF/svcMZEzjZTXx6tMha0x/ERJGU39MMBy/wcAVjDtWrYzu
rhyT0vLaQJmzmRCYYPBXXWV/Ip5equ175zeGKbo4T3jIgmO0LtY3OCXz7FNmPmnWhI090w5bjaHp
mciTk9aANs3ZYY/stkGdse3VUaZmuByd+JtgnejwS2JdINW/K1fuw8ncWVjaAz5G0DcjBQU4sp7N
f0UqbGrtNvYq6YDVLmqJJTaXSj05bnA9mO3HCPnHPcf5XTNPKb/0l6VXhiL1ly5FnAKifOIi0ywn
evpWrZrRyVt13JQp7gAnCjVd29wjDqRukvvuXtR+cYqvZgT8wuaIflf2kKioJ+lvyKnCYdKJdu1I
ZLUFjVQKviFZyE/qTQYPElPJE9bmuVSATdPnBRR0T1i0Hh99rHCxiqKj/iyZHpcCyMoDchU2GuER
ER5di0mHWVPe/xD/4LAQIUo9dKOavWHrX4Est1+CtXi6JUxlGokAGjP+5MIBJO39hGahKtS0jiaI
BMFMJASYKH6yi97dfGdIILk6W2g8reNHm6HERkogc7LO9NbDfFlKnUHBhU7B2+OATI8IcZmEJSy6
gqjifDfj0XUNq0HLyjgOByyxbrUxrS8LBcdSyYJvUo7mxXsIPpgnGj7VVxDGPhqZfHrieyWEVF/R
IeA4SqvKVIj9toLe59QPFM4VheClJOKNL1vGFfZp9KCcM/cihdINLoOhTd28xbAtPFfPxe+h6yri
/UAFel05H2Cp9pyS6G+YquV+atjRwn+VHiPag12Fgy8lJdcLUQLXVDcoOOxTgU4R57NMnbpe1tx/
kzrLXvb4PE6NJDjNJ/Mmk8fXz44xH06e9HuFhqtGhBBFAsXOQ1yh9iVTOBJqarMajn7NYbt7gDoh
0Go8oT/W0RQuItchALAfzbJYhNyxRfQzQeLhIsH55w1z8SUlwsGyECxJWujbrycev6U82BlQrU2D
qpRrSSeWmnFFYQvbvZwO6Xbay+ogo477OQ7k54koiEw8QIrw98qA1pkX0SkM5Do6MA5SDP/dW/mP
SyV+Clh5D1Nr9GCl0mJhVirveVljDsOOH9XGQ//9Uoflg9JzcrNPuBhs60n1qxZF25bG/Lkb0qFv
1oopH3kiD85xFPTm8pT7DD4C3V1WLXy6KvjMpjmxauiL/4J+tNhRY0KlmRrCrejkUpotCAcjlRw7
+9Nw30rcm596ZoX/DyeKFEYDDLeWq9GOEY79K9NQWZm0Rm37Xecmp/2gG9sC+T4I+erXGgOUxOEf
gKWICLpaLAnbltce454JQvj4H955ZLkLRNco7DVH8NH0fGXdbKfplV1hAakcirnqWsFuSZVOEA+C
QtF4tpvINzUHUboaCVXTcbklk6SO/FR071mEtI+hIYXh40xIgKRItFFGxkX+L9vddXztmUpuCasQ
CK7svAISxIO/Td3QJCBrUYGyK9Kv24svYWg56RCjThO1reSDV/8AA7RtAdUqSvduiMW7D/0gwP/U
Nl7yciX6Wr6X8ZWSQnuqlR8eX6rUUMAGyxmoA0UMynvKHwrO1shjvI22Dva1Y1ktJ4KJzfuZ998J
cMjyuKWZyZiopPBm4p4pbhwMRPXI5xdlBUzHkSJs1HT6Ew9vIInKihPf24uzkmbRLROZEICscqGa
RFPnTxdIf/xoe4cdpiOr02eU3VN7WNfLS8KZjX+GFlNZiXoFqRhOQAhLeUpQ14oGarvHKhqdnFKk
5ZPJHOTTxjJ5mH0CCaRkZAEo/WD8JEUTGRtRBuWnzT2H2JnY2sTbcOgdtRCLeu/rEEz4UIiHVdaU
IDP1y3vR2BJ/HABjaTOq20A80Iw9CCKtiQUX7jp/UDXgMD/RUl0xD6D1CQkz4GEhCYQ/V0FaeOwf
0QTZ1/U0MgGkEVi/cJzB2aQ1YvH8H5OYrUxVmiSveaPZMSaRvdkUS72CHTjr8wT2zLufIcnikSbk
ufeH3SjdBWMp82/aEw25UDnEdvc9ViROo6rQ8KQc9DVlYU0lrVS1cHCMNdEuZruagWIZjxSaXxzp
ZQRyncKoMB6Jw8i2y/7Ku94J49XdgJCAPuTQgQW0/TgNdjJkoZu7/5if2XqbYwbRxnL/wz1at+Rz
b45BmEa651HzmAteDEA9UZv8V0CV9pY87IWVIoNHNO14XQXtXIniZEgGp91lcnKQKV4MhNflF9SH
fUdWB0vbF5iWHo/HlsafWGRdIBb4u6H9x5B1vkdSAi23iv52iAEpt9Q1fVUiH6MKuO4k+AV/egx7
BCko8mk4hDlrRyCpMXdRZ00/YcVmMY/DXOzS1wUfo2chvdL/r02KOHB1O2F8s3ryQdnzVkFzsJ1N
c6S4f//3NDkJqc8gRwjEyodk5KfNZ76M02H5+WylFfuJuF47/5+k1c6ZBg1xfzXmVqa984NHjMGy
tpwNHs/O283OhHxKqWsYlN2OD40Q4rjD/jocsN3z/XkDzOBvHxMu4GJcboRK3Rd4SplrpX5poB5f
7+BO3MBUk/F65/NmiBOr9Wh+spkrMUKLBDPn6G+KJjE3sgAYqs9pH5NhVMAu2jwkzV46DmUidMeg
FPbPyiz0CmdiEeZ/OOi3KdkrocDqs+LsL8kjXdV3/6IWcLGDHNujHN8d0JIUnvaMm6WzKtuvPF/A
Kqh0qVEOEzOQSJF8og7JF7N0tZE9PTCTbrSjztmQwT4zMvHrj7bEY6YZxFTUd9LLxOPcP/YBzAFQ
taq9Ah6dM6dZ04QXfbLcliD+FESGXh7N7edI7eT87QZLOOWkZ9uoNH1Hpyy4P1fJvHWhhdLGPpn9
6bU2qjwJpWRIvpVVCtP1WHoj3EYfgtdu7Wt9OFW0RPy4b59dmG+mUalD76t37vRw4VZvcbzZGKNV
nmzQr8S9dBXiCu6SjKNN+7varsg77O1ucBzxSu45yvB+EbKC2HIHWfxs6LWnwf542MHgkTRa6rvi
Exn+i/DFiKenUXeJWtNWU7e4Ky4SdtHIS2q4nR5MtAO7RE4NPjxmoBKY2cS/McAFIRJY00sQIAeU
vtSU6Fbspte/5mYPAJc6hE4KWBThz+Q2xGw8+ncqYj0nqm9xN/aCngxOEmNA6sxvLx5w09eUsHp2
BqhsPphngHh6D+NpKimoRj82VryMLtNuchyu7RS6Emm/kKsDpzzSjkdR9K4BNYnJsdj9gIh7L5hl
5YOtqKfhz/mHgS7by4eEabgmOFn4g2YNmD4HWC4CB9DyQXy8Apud1wY5iMbEpnVOnoQM47JEvWmQ
2lZLGHXcOc15PnPriDz03inEsNWU27e7+Z+WJ6THIPtAAVC4M65xyAL6L03AdwTKXTx/wHgnRhOT
ILE6Vrh0xCBPZmSrql0uWMwI2UcBfAddOkk8QotokrFZJOQaIKWcmtQgPYhDCuZiM/bAiFgJOq2L
lmXCeQqpxwzmg1cYbW6L5vQasqsFunH7376UYWgnjQSDV8Bob5C7IW5J3kT8HiDKXlBWvtN+83vM
RXUyfqKQlwzIV0QLverYE2o46kjkHqSXoni4CGKUjV5RjqGgjkEVW07cvw3J6v7k5VsSEJAVUirE
8GvLTLUui/ayHCWNfFFBqMnVKkuBTxuLnnNC3IX4c/RkL3d4SD5KIjQuyu4gkSvEI4frzkHy69xG
BhQ70uSQwLp/RnLk+uuhToeCUW84iO/Q9aHEurK3NQBaWE79MqHNBgJyee5HjfiVWshBW4bCG00G
sN/MtNwOMPFT4Kt8MHxefnhVH2qzNgq86oaF/xQLi3PX994KiazoJG6fgtmid6DGWjI6vqlDfDR7
wapEgtM60FTYyfO+t7ZrsuWu7r540oHMcu02aBhHOypAwiWBLDtXxYc4guIMFKoPsNDk4SsP2Qy4
oCVVenNxQB3PlAVsR80onX9ZaD1yxpUgieOOsfNmgbSRsHm4RFWTTA4wfJz8wIjpqZe0YVBgqNPs
1QmBlMQwtC7kI2KjqG2PgFPmXM7TKA1iKQfSMH5RK1NugHQIBFcavsBSqi2Z9f9UaucaydGaWljK
FpT7ZEtOkzStj6TJC1ost3Xl5jht4S3Kk+tb1cgaukiarOvvAciUCCTQAdXWu6vu8BZn+0XYnvSU
pTgM8rofw/PnzRlKa2ZLXOp/5u9aoqIvGMM5nDWAVQvHfXrcbE+sp4PMWwJfpx+lQM5jASOcFuIp
1qqDh+PD541hM3xUlvoFuEw+q4LQSfdUxp2MOO6rmVKlzCwzl6+3q8yUdYBH+Wyp7U0iT1SRmbre
ON+HWrdIbTINoQaWwnUjnKrMkwmfcngOmh73Glh6OH+yatRvM0FAqEYJ8987/v+9D2D3R/ed0Gn9
PYcJkReD1bXRykvddccNBWYqm7gA+NPortZ8XcapZWtojqFQIQmCHka0MGHHz33rcqDGZz0O8rJ2
Pdm9wnLEddnn9I/NQmvk32RWA3pTjSUJtBE3DYj8H/qobz5Dko0yI+jClpn4OErw7cirkJX9zxa6
oY64DITm8nBFPNKXkEkG95n36tawkFlQ2Te//pghePtXkeUy9B6yNSGZM3mPIzd7gJKogBaqW8OX
LzTiIeeeeuCuGfAQvoHMpyuebX1UgsK4HwE4IDOGr8cvaxMMbEVOCrrKyuBHzegsZqrzhXfCQfK/
CIqR2sXwNgspWgr7qAiFd3z6jwRzuhT9laMuMXOMPEHrstxAezwnAx0RBqxVUI28B8drVx7nshg/
k0twgRZY9dGQovxRpOfCWkf9c8WYJYcZyG658kuwURCJNPCWh86vzJQYtQJSqJHI/Czl8J2ROEBF
cBbMRqsA37nwZO5j/OOkw6n4MT4cr6NGEPfBKkqwoTTWUhvTnb9yTyOHZu67E+CWoDQoIQS6Mc2Y
+4HU+kVBVenOaNxFnZZ0RNle9GsKY9cHOiVGdRrkxExjQcPay5LnHqp2fU7M6DlA8UzCsVgJSLE9
yJQ09dHxIdNqxEQpL6erQeai1tFoaENhufR9lPDs1XUpx7QUcZVTiSx1Pvf7a02gwCdf/Ne/xzxm
i1eGYAXW2FuNrlIBxXz19SH4vL2dmvYwIx7p7qM2KjT6ali3TSRHjrD5z5EKua1rf6ByG+lPA0gi
EnJCuxxFQRSRAygZpe9kHFqM5wDloBQFMKNPRzLsGEgFicJRPJ2xesowWis1zNmHjavZ9av5qhyY
QJTB4A686GHESLdNzpUIZPq3DpG6+FNckaNAhUHCbLsDp3mZ4NJWVoRUDEfGgxn5XRz2aSgB0JAo
3DPyD8tbstCL0t+4trBOlW7YiucMKTK2hDzdXV+3T41pGgPPBcqfnpFJfjJ0EMmbrr7FOImbWIsX
4tm7OvX1GNle7vEFS7+D93KbEJpTFG1VQy8CnH4RU2T746ID1+2SZm4pPXfPobUpfMP60dhnguh4
lIdSPYThJJ1LDDQfl/8O5+BBZdClzD9Y/OmRrgKqEOzpQbs0j5J2aP6mBaQVXkNqzDFldjZect9I
9Npdx9iT67U3NXIJ45cggnfWSAVpPeu4A269quPoEqnRN3MthwZKqEG4WRCij0gUp6cVuLrf5gJG
liokOByWWGBW8VFidoIAgQIpaXmk97jHLImdtwUnadywNgpZroPqMvBnqTmeZIgL9K60YZLwKve7
hGZNzzuU+P/iXeVBPW6uGqqnJJtiEd3GZpkfn40GS4MmBLenNGXN9JaqyKBp9Ll25L8N0jL+mbsR
W6i9isxD/0+TPNP0ER9ZTXSBcxXCc9CTlHfYiuE/va3a8dyT9UBxqWUPqXuMhPD0hJdt90//wGWL
e8dv79ZADsUN7B8rqu6Sfi2xJDEBiFTtAVqCjzXg1VVvqNbuLry6nUCRtTk4dwteXPOcp755ARrL
vsyjXUM5nRLbsjdn7lOtuEAPOfCfXpwC9jaL0rTsE3QdMxINKGjRNAcvkGLEg0imIgUIeDlwd5A7
J1De0eTgXejshzPQy9AUN7WcUdMRT7mD79fC8mnRVRcY4D3umLQu6SaJputKZhBZyg6aEqE0gDTh
avRrA3jZl5ELacD4L1MuvweNfBkvzHaQMTHaYu+exzpn4KntKnAo13+6wPUOCVYSpxZBClJHRA6+
fZfuOYXyhbMNKY7jjZoOWM7VFxmhisMRJmdnz8UcfYnjvd1iYci0HtjX8h/jpSOdAyLJaFWQFlkE
ILssxfZFOy/dBw+XX1CcAgq5NGY7vHd6PPBipMvxbkQ4nKzmhza73mXDeDqPRa5PpWKzUSbwH5bO
6VvAJwPrZOaftztzUnMYfYyZiVuxuKiYcIIVHL5KKGmzP+GgSTPLbr6CsyGFuJGiWnSWIL/4DHbU
BheNRMdyb5wCvWkhoQ3bhvT/bhn0fn533GOJhoLwVS9eAdYkWd/v798s9+vFC7atXMvtqAePVeIh
3IdacRs8fU32pR23Dg1pwRv3UI3yt+aFwzl6YM1Wz4a3ZwT2s4ldmTrY7MEKY/wEoTrs/ftHrP77
Ttd/y5b9XU9tfkh/npEAU2A098OrLf36UDTFVL/7+op5BqVUYhC3a2/GRMSte/zOkJE2xffoRT0d
GZR6grdVJO5EdfQk4wjnAtMQh8DQjc1a260+LtHhCHJ/WIxpPpPTIsVhRl4GKyOf1+8bwFfdyUZI
nqcH8icIM1i4YmPvhc0Ihyo6GVekBiEhIGAqoZTrtP6JGVuIYqiwIkxbb9d0RRWAWe66AWvVyabU
FJVWpDcosJF+p6lrgUh/KNdq//s+oFEXxOEjlc3E1Gq/ko6qhMCpSIsbUalvsUJlIHy6bQ40IGrd
9slikiibtbpVH/3TRx1loUEUfhcdxp9gH9PEWN6xaXxJ1WWdBAbVahLBBJHNNszjdX7O9WG25QF4
sjjhpIJdpex70Fjtn+dC3yfRoj/sCr2JOSO0Hy36A6dI3iXvRdJ9z3gKaTAbO7FdUWJHl3x9dYMv
zCCuOfaCGMMWpZfcPKjxIAqMyNvioR9lfKvtTpDyjtL/e2/F8+MpyoZzSeb9RBWG9BuUwV33DBiA
iiKXYKygTp686rqWigvcAXcm5dbTJeZ0nLWaiT6zlJWN+3LBcipLH0ZKiqFt0GBT1MFszB6H9jHU
JbNLrje3hDUeMLzmCOsWM0TVPY/yL++20oPWmd7wrmwGU7g/56SxiQGk3xOQFkTZhLkLC27CxHPE
yAseFrZIS19HxYJqs0iXgRvdoEYICet6vPy9JusNGpHJC41gYxvbF5I8RU5Ur9CzUVMPPOc16pQa
DG93yRMLh5otNjMivH+kuiUzDJ10JNB+rcEgLt0299CQjaX2QV5SNxG69eCED3MLIkTuzaOrwqkn
O2HKO2LMFdcvv4od1a2yRyaxUsm9vTei7QogyaQXcKeWxj9dffcQEvfUezGd6QpF/SRds2qval/n
I2YhhBbmpCWyZ/TMePADoSwlozuumTYCurmN1XGoUCUqHF4qLbwDasRDVuUzL3aXwvqt7uAMqcge
FHc/ElPPn1a5Ws4jl97R4WFXD1CI+zU4CwdWG3tknrZ0dOOCBZQxrI5woaRoqMjxnhB+yhz3XHak
+F9QQGB7sTOCgGkJddYd9J1PSBqLT+HK8dGtVG/yICrP+ErzDlKhrYm5RFfDFtcBOTJSb4RS05m4
+Wr4OqD5zgYFVnp6uEOpUCCgP1Sl13xErQwyJ3IK/N4b/cnpinAzjOoeCq2XPdbwEmIlPB1vzuSw
MJ45o8V0NMU4x5XgoOhXP0JdttFExnJpItw9G+OguUcR3Mf7xMdImk2Mwy/gHkA9Amb8aF22860j
PKpWG850q8c6JZbLKw4e4EWvScQ7rYzyLqTqIaKu70GyScgAHCoL4LwwueMaQcPNVU5gXb5N8XWj
poNxCTSG4XDGyJ4pi9S1TCZslPV5bsa1C1F6gNaeBc8k/W/3/Q7g7LjtX9yt8OKh0ok+RBXPci/+
cpuqHc2cVYLc5nTZAgEYwtbQ9i4FgaXBg9y1EoMlBmlEM6OfqFIFy6L7AhSUyYZzFxmHvgMjqGZu
qvTlgveWbpl3wfHySyN/Wgq2X+w8snesRVcHcVBqdHoxdiqJYCjQY0p0L+Ue0W+rqvgXpDtqrJ6l
rlse55y1qbxcy4bCdcEFL7ezdUue9NxrOJ4a14vM5u4E7iyjoJYS3X4X+WBQ1Gr6AXt6SP6AeyQW
y3gbRWuqcaAnYk/E6thbHOmI8u/+E9NfPzXu8a5ajjOCBtfU6dOCzfLvVvRnLOPPle1QY2zrOM2+
t2bv7XzdJuJuFxif4ZZlECL5CNAkQJ4awWfoh2HxYB5zHvYGl25lGkslS8V3NoRuu4svu6U5OlBQ
lHwqEZHmWZMwXc3tzLQ078VyPs+o6Sb9jhwexj16fCFqwQAxk2MyvNCqivJTbzUl2KMbRqywQ0SM
Gj4k8yCOu890x1DAs6y7cYEi0cF4CjbyqKmY7I5cfjwmmF4/MBpzCFhaUPNgq7vfpCR0e1Y6LKhM
SA/RgCNz21BuahR2Di/Hf0FZppcPpaCEgTbmdsWt4fqAvrTCtrLgHm7zTnNssGYvUdC7AemOwOhX
jnybGhajiyo99lfbgFIDljQ82Bz/ZcCedIZ5jzpQjacnQXKPXiwcIjTgS562YpwCEzTfCGA+WUGh
gB7Jq8J6cpgvHTfpJKNcSiYOuuSsSykCPAGwZV8zGfD5Q1KDmsEs4jCyuat0RIpLNG3baAOaMBhX
CMekRjOGmyUsuIoCyH8Ez8fP7EXxUy+7os2RbvVVG6/prvnS05PIdWGr9cDHdBOQHCC3JSEbb7L5
i6N+4busYvPH5OfXlCIDPocKlAPiKSU3wI91MGP59u55QphC1fkEp2DUNmX6aWlVu8FocIhQlJM4
ppwuusrjoEtKLxwWGYW+5Q2ZYl9IPdKRJXOjSP5CAyBf0TF0ZsURQCbyWufAvzuJqnWrbjlvGAvn
yPDOZSOCdoG4bbOeAFOrkE8PpnoQm4AnOFazmdFb7z/G/GNgudrGlWaCT23DvjzYRbQ+G+pMm6nH
TjVysLGVa9nqYoFdG9lpeyopZqMH0/kD4PG9ROokw/vFfc6QJg8s+Ntpjvqm0GAAVYskEzinyTcP
LaIf3brypwEh8DEVBDCsBQnK3sF8sFzoKB78qi1uaA44ZranVCqb50NZxtFcujZGsZrvTLeRho8o
baaVpeK+y8Slcvxe/oHRhw0TLdIJR1dqG5XwANkroU+Ero2uZ05QKh7zW+ECYL5023KXNXoht139
POo8o9nfuQ2jZyj5SOoIh+FgP0mYmtHWcAstvTxgqNgd03OFwU1I2aTMYIPX17OSTZTFIGTm5KMi
HmAU5CLxlzKuQBtMV/a5I1znSQKCAK9yFdvr9q1wAs1DQxLgPeWPN0HeQZ4XLpdB6k3uK98pj2e5
xExvaXH3KdqydhRrc+X+VvCDpsu4hOubRZvE1i0K9JXdr+w/M1eOq8z7na5ktOitmi+UoRJMnPoB
h3xloeOeLU0t1WWS2W97B4GPLSDTp1R+UT59vuAp7lj0eFkWbG/izh6e24DXPhupDmiyngRIq+Z3
q262yPEH1SiD31eF3C7dKrwOwFQrvWcerh6YOJa6hXMeCgL8/zxoQJkHGNhTrx8aBVayagn3iA5p
XTtk4NEDKXTDmhk02Pi+THDp7LBccFvq39GHtLc1bm/fT1Dm7oy2uSdzOMJnXjnQk42o9fkBAtRS
qSwG6nlef9Po4TTRnlgDddVPbucPf5Bzun4boE5ggyBnR3RwgYCkH6K3fe8sDPx6zsdPeevW9wnA
GysmPfU3t10ntFiVGnu/9O+PaXwy9+efJi2yR1PdRN+AoH6BdgHsUYizF2qlaIMGpYcU6pWiwb5C
jnLIwRxTNvu40XQuePLmxE6889WFuJUZSAXh+mEHG4gWiqU1l09Uz2u6Z4XCF8H2mFnWR79CgV3X
+vD1H46TM+ylJvM1/bmsygtV+MCzi+uZhwJ5b3DszJO90v91yhAaxEM+V+2p+NUA6x07o8r9mZds
fRl9+x9MO0sxAKkWgMDeMJ0CB2dK4Fwkdt7JlxUMsvRenlTeKflAlQ1hJMXwV1Y/oZdIcdmoJYPt
KCN/gi47czRDpsBFYAEvzcLnCYQbN4vZKnIC/RVF7Bj1rxPN4SbyIlEzsYZDMl/tu0cCk91LMxIb
T8MXx7fOHAhIb9NBpksXHIuC/3SSqjUGM7a5Of9UJM7pZoItUAiKC/EuIXxNX3xMjiAFdFygpj5l
1puQsxhPNMqKZ8aYIaMUubC+pYU6uurySmx69k9FaxF4pp2A02bAmVqfoeFwoGogifB1SHdyzr0+
ew24NfexFH1vnww7o+g2sbTg7eZ8UT5v6jzK2cY7/5niaVm4iJWTPbDSrhryTZaykkTRDfaBLT+5
okzO3WeGtDd2EMwEeXor4MFXK6b4w6CVpfIr8+kmS4rbuT79f/GOnR6Eg4JKsod3W7GpHLLPbtj3
uPoVCemLwkX/YeWv8c0ZJbC1t1R0LiWbyh3K8XeTmZESDoYOTmvkrNy51ceiGBYIr7XHAygDIyBP
ygeWL0y2+eDNUAREB+V2EIUR5w4rzyJrF8m5nnrgIFixGnEKnYAKntPLgXbBLEGjj3TcrKcomYOf
FhkGpcCcYn/+hcprtXHxvzRtSFeqNoo3QFHtABWkSFdP3w2gQ1vElgciI8fzrKvlAZ+Oe/Y8+b3U
j7Uf7KA5D/LEDsmWhbwl5nhPbJR59ALhFGfhlBTbpfR3M5EVK2Y+SKgJilWEOT0oW2nRWvJv8ctG
iKdTs/xz4LdJxamate0CM4P0NtcxNSw9FbHtdAi36Y5srtBpy1TTS2xhxkUsitOaBVOPKQ05YIGG
UbjWwHAqiI/KsFpON4AXHOYALpHzBEeF2uOAuNLgF5CjPqnGvrV9FeZvpBQEajrJ0ROGx4jOO0kf
hrr7YD11ls8/ywMEGplgyJsHaThO0H6jS5r0X6qYso4UhCr9hWxRVUniWXdN4lOcwZUvvBSgVMiH
23rAzbjiunMvban6ZzW3NO7kuymUTNv6sB57b6HF7BFxwQQYVrYxcqFb94PluVUG8Fh85mdKgEYx
x8WpHqxm1hmdPcCOnPvHWTGMgUY00LdscAeukpHEH5BimxBOmN3ws/l4WEI+2vMUm7v2d3Js/kaX
J5U7vI1S0P0L9ZJXPbCl467cmiKYuOV2RezOdua3r/DKYsb6UB8a96H+BKticIbq3LwZOuJJ6f0O
eRCDaVDTDaFy9F/ohA56sdOgDY4XORqbP+sGeQcpOZxeym9mnBJc7zICC8VzURX8mdIDlKjgTR7b
kDy9eUSd/QGkBAL8Gg5d3qhV2VKWVzTUZPlyDpvBcm+ae6oi55Goh1pJz4au8WrhsYoDZw2NwjFn
1K5s02YgxUd8ox+9phpBZEql3cR8wZZbQaJyAiZRSENFcyjqcWRxGfyXXNhrQRzIWElv5Fr9HVS/
0nlKCHatdMO98DzSAG9kIftEeeCi+H+hgSh3b1a7L/YUAz5KYN2+vpnoctjkjSftdzlN62aoUuu3
J3TurqvyH0x/HRIc1p8voQ1HR93B80GiG2QaSCToFKqqhMDcg6z5Y+vBsHXb3YMhHoMHP3tPTEyd
CPHTJdUAFMFJ0V+pvXVj3Chryr3HkDtoo957AZh11snkL+w9pRjd/XStaE3qrV3IexuyzeJqSFqz
IfOgk4cb4mebKAoe/0UHCqkFO5yaSyxrcFaMji/On3XdspEyYoYs7GrMwJslF0QkhLFj+hMLaEdz
9vruFpQGRrbjva4FnLtYriX567tC9HnOyRXJXMz9aA5MMYYdOINJtuggJeZGOCMQG2MJ3S/7ZZZL
95sF/TvoilUV17gXLkRIP9jip5OBFfY4I032DuOhRtzBaJT+lw85btg+KU3xLIHe3BXP5F34/+as
sddR24rZf7yU8PXu3YHryUvApEvSQFS3G2SN+edoo3ixiFknrgotcMBEcoof0AjbJVPWPhmxcS19
RrpNLesg99ap2hMTT4y6Csr1YbEEZoD5ZljS8AXXVnwx1OilxjRIKAXLrUZDtA7ks2F8Fzoo0+we
p0GXqvjLIMTY7MG2QQNGTZkCfDstmzCibk4qtfdeAZ5+urpwdh5V5fVkqDwro2OOmDLl3OPlFc2c
uNJCd+JqIhsl9oo7619MlqcOB+tb5lGZez1IvqI4uedoY/7G+03xCqH4rht4KCMJnzIpRwT1++VO
UkwIuY+G0Sk9Qs2dyVNsMVN2qlw3co3c4Dno2R0a8H6L6I6x9ipYiXSQZOBuJlEbvhIearRF2/Oj
NucB7LYBwpKoRv4i13oHlwPl0R0II72MW9uqXKcz5z1Tv7HUYL75+UT2qfu5JZbylIMdHQ/cFO0g
MpiKDHRx111i+3pL9wzcd9Svaem86DpTeBx3jUhIU+BBHwLD/mZL+WGLeFEOxEWBDlBzshBaE+X9
ZGWXTgZ6cE139wafw4XJIJ9tiYAP+xyhRKLTyYwsfZ80P15X73+EErVaMjuL8uDDPTZ6yVC8pxCk
Lhsexu2du4U+bAPLN2rccpY1lR96PMUoNDA8MemAOYMbw0MtAoTTTrK9Vq6RuI4w2ErqEeUwlaVi
N4EVPXUIjHIiM5W0NieUxvW3u3gGIsS3FarGyw1DAYhc6D5aOfEfLqEwYftge3mx4brgGKYJ4d1q
JA5vNF3MMKBr8BxlhT0Spu47d8vgNWUUUeKJ9+kZbv3Vhyq9J5xscV9S1y2OWpyGhz3kmd/y7Pn1
SneDc0E8dSDHuIRmSd+CV4Zof0+E5eD78W6R31jLUIlxOH31Q25vrHid4uMhDGgBZgrDwFKy+2P6
/WUT86oktsl/zeBCzKZEeaXQ4d9pyGFKiT7e75/yMSNu4jhB6Rq71YsTM/Crrj1zPD+ZxXbAPg22
1Vno+gYX8Dsf9aKIlDdJ7GEqZk8xiVmTputpvr0OTp5mlKgMACHsJPMZiquq3JCuZQsoaFhlsdq8
lReDo2yR7MxTDYz81AVPVnUouWVPBuRd3OpOnHvq1TY0002Ilyc2Da1sSEoTHHD2jJ2QIQSuv3/X
ZNwgW52qd400iOUyP5JqjTbAc1dnCP49fKTiKl56P9bsddAIZke6d6C12NK0oa8+oxzkcnAFplJ5
tu3kcA/2xEOcsT+56CoHtMKKk9isPGKJSviB77vSh4bkniPZNe6iph3RuTfGnkk92A379aIMp28f
HNVnJurXa4usI9sJ8R+R5WUze7y6D3IdZmhMpzpfn6nollfcNu0hKLLPMm9BSS0CMRs6ipkR3XnT
iMHv4p8vyWRSv5GKcMLL1/xe4Uw0Wr79rx/eeURWNc9A23DpZB+8Rbw2YHtxP1BO/5sOZqAz+3I6
dtHdm/rjwrdUiGRopscOkwaZoUG8d64uLk90G44cEGPOC9ANKwXM31HLZ6X+r1GmgX7nmhEbN/WY
lX9tTzdTMRP88OKiOZAv9O0szCHwU8ovP6jXqDA3Oe46eqVL3cRvbLLzccENOP/narBZr/NVtv3B
GQUrVb68i4bimbEu0YgG3Qh6gE0AWZS8yYnooMqJe/pzGKg08MnXCqSVf8WUKCiMF1N8jz/oJ0HT
lIvCWUV0ZkhFz4IhHmMQz8bQA2nI+Gr7A2CccAjS84xyoaKy4dopPvhs+DT8P09YwYTVKsrHT2aM
z60/XsiNxV9IEMmBQ47vN0zs85EkDNbDxuEQDu5mRLWGiQSIfZyfTHjUsihYHa8YzO0HrDp4gRw3
YCCKjtxUI1i86iZMEruKAS+73xDkBmOBOc/9J9XyurYCqeTFKsEVT9SPnYNJ+7QAabEay5Hme1Gs
HmQ3NjBD1ujYcIxQz3QT+rC5om9yGEq83/A0iUn0iFvmy802GeKjI1YlS96m8yJtfxa+Y+Jsr1oA
VTaM6YoDJc5JPhbosW67KklHgqjfs5ng2VMbaNdFwATfWEXvRrNqN6c3USyTbMWTUU1RHHvExpCQ
B/faBMDD7tXVZ2FiI6QkmvftDwGUhoakwrhJAEG6OcginfjWETv9YDLyVev3JuprlP8RfVx2xjKc
3tY+pT+EWjAbEMwgiOcV2A9x9lI1ZyJwEzpEMDA2/unSsLxc85BeAFnQgc7zSRmggJ/UJ3UWqpLR
QxwifzeNEbpB5XWyCOtsEZ3QocMoi+3bS8InRlqeBQoM6fAeCV5sc+jLajAOygjQ1CNsCn5NXkEf
NQE8fH2VL4CwVfvmlxlfA21XXWdKTCKOH8RDdi/1HRUIUj8PKAecG9UYMThMsAUm0vJBZQup2mca
hRUBMpSe12shqrmQdPC59MCL0ZE8MRBmZWgd52HD0UsKdm8IPzXm1zLbV0zsSPr3qZGDafi5E8qJ
W7E3EIKkQRpuEm5or4zty9HMLXZaJCsfV3VIixJ71yPyPZ54V5fvxPgT5a5Ee2Suv+Uh6gfrs+T6
Qrc6uuLwiPfUrNdrWTCvCDRQJeMDF01lNzjkodHaVpXEOOkgeLuX/QtDvhXVeZICLOMAj86aTwuq
YPZGW/hcLRhuZU3pQnYgogQUHrbfzH/60nTl3m8ZPcKDK0og7Ef2p4WAnTPOo4wRr2W/5dGmsZmb
H9OlxNfstEUS2EYaFGKn45xXJVpLf9D1zQPEOcJ3ucYPFYnHve5j/Mtdf+Agsn82r1EiN9yxMMxl
QfkPDtK+b1c5V2lJ6MkZ/XUfMuh1AIjCzvV0lj1hi1gdUrVTf+hXO7XQPXQUOdMD0ToHLsC6P3mw
hu0zdHeHpzzlyXevGCZ5NAJrYhOGuVM1iOjfNdxVqenp0VV9olm5lIk74b+EtY/oIaoJoQ/WKcqm
0Y0c0X19Fkz4O6Vmni0YQZ7kSdv0ZKcEWKNiEngiJMW/Zi/HOy0LEmdrBAGM2IPa384WLdwMBhu6
hzu0sHr7Fa6zMzhPXFWKvUAu5f1cw9reDl4Ux+DiLkSP+Fkl7c1Lhq0MGrgeE4+Cvnq7t/Pce5s0
c7D5Mkoideew262c3lVtUZfjBnwnbRc7EIFqrBFdC6XB5x/x+P43vw1q5fV7N/011kwHNZhJP4wn
MF3+57H02pUR6tlWDgPs1YGjrkXTjdRu7WNE8cTLKCGAOpAGmO0Z3+Xy0CbB7jZG92GsLdg76BRJ
O0B8Ky3UnyosVd1bBmGb1KxZ5Zh9JQsU5LSlpX9DVWJsnnj1DBMHiUFUNHg3sJaz6HWnAJv8cGcP
1p6qslcP1LwlKtWpmGy/JkcHesfDN+9C5jd+9MiwKfDFLG8IFquvGwr4UT64AR9eY0eu1h5CVGGv
MtjA8j/2UY9olVh4pkUc5slS2Laz734E6VL1TJrca0dLYIHCFb51L3uTxFkWj8GgdKRhG9Z8/kdi
14WxtHNgEPWPdkkYkIjUVVnUKInBYaOgvKnnpyJn/r0kgCVCn7CIZUu9MWINOS8oTJaRNBkdGbtC
vTCXDbGlZ7btz5qdC5UZXznioKG+3GKi1c/KyeqtZXdnnIkFvs0D4S/e1Bg3KbzlROIGlOdP7lzg
5axKIG/Cu3c4xsT/17d99IZDkyV6MXqX5yt+c+aUiNes5o/EJQMlqt1mB0j0tmtPiY4eMnV9Ypsw
wV5PYuhLqwSH75X5nWPWm2SrvdZ6Xdu3sKwki/EY8uFnOlkfZLUzeRZrFlbblaZRjhS3CdT6jI1L
ZZMLLAwQUeGIjNCZpd1nbvNeuHb7I87fqYWA7/YZlOhypo8lyU06BPF97GV2m+dD3bD5WcIzwPLK
qvq7sUlSWLmteAN4YFB5zr1J2lwDoV3mZoUf7gjwixDg0ge9kMnl+MLt0aAyYsdmscauwH8VYhk4
7NQDW+2KrWDyT9QyKUywcEDg6bITD40Az1sL1J7pqvQyOQwypNqKOit42OzL0Qb4HoJLYempgnKF
2OTzP9K3rTwbNV7pSg5FQuRuA5wg2L+lRKKsSoPURhgeLA9l/L67WmL2uFyxWsPUjqOG6xC5qLB1
X/Z2YvBh9ZHPeXmKUm4VZM3ViONDmB2JCu9m6uNMRj6Z3zUSzc9EdRJnUz/zGxFYxLNsaGRR0ads
fzx/G3Yoz52HjtRzzd4FpioLZoqdjMTmRXNG9wfQk81oRzo24lLhYe9kEIdO7oG9S01EFp6N9SqF
Zx1++jgE1WHuLODRdfvivxJ3L+LYlg+P1kaYFVZ13Wz+QV7BK1uwttiVSGvLu20/QiUwDLVGRlOK
A8y1UH7+yE2to2pdiAcKIYfCiMrDM+ocqSzyni9FnOu8+4lyhqlN2P1opQxULHloYPzGEYfYK6HZ
8E0iv5U4BmHhLia39+0Iq3NHrMevTCchHPxchlhKVs5owcubPGhir61xcwC2vpO8+Lfc85pr4xZX
mzV9gq3I6Q7qQ7/hPx03693cB0bMNj+CVMj/XJ7i6gMy44EhyE9xXCfgry2Ij5iUjpP36Vs9cNSb
OyFacl0nUV3layBCCMR8NTqojycZbNjAeh3/iMx0Z5rYCX3hA/tsVr7XE8H5HjEnDy2YXOCtOdNs
Tg45eNMSXbsYAjlZWpr6LZ4FTszS+zvMmUc0PC4jPGHYEC28xliIq9h+WHy7Wr63sHt8nI4ByvQT
EurBlD0dUUNmHgGHfkg1a900CZidQ4MQYCphmoOjLEm4VFhnNy9SeJx3nzPROh6ZtCZ7Ex+EYE6C
fJhd+8pePgLQ4thbJ7x5RgyM3bCy5E6+uTIWPSrJOWcs5FDpVwyxi0hhdb23Ak/kWRQQm8YDsC3V
U/JrW24H6xCOzfwJ0WzIxTdi5Jv5VGk/M6wqWbsFG5LrdjaPCGqT5JhHU7duIvM1d6MEa4/XLpA7
qZHjMdshuuAMJhuvkYAxUoPhT9pvEPVOQMDpn//ZQQ+FS9lwrtLFTqZlS1/znZwsoy8MT82iDWH9
JaOtikS4oamhSkjEoZ9riaqcyHE1wX9rcQ1YH+pnyjqVd1GSCgscELgMG7oeApiL0g9Sz/0w4nHj
j7zuR8yTJfUt8TCfG0hk6qZfl90X7DKl2tzk6/9mCBH0LESvCSaJgA6h0c3S9UQl/9TtGr40/EeT
gQMWNPcbmFonsbWashqlVUnodjriuSsSIC3X4xdDdgZXrz8++Vud4GWUT4kwKYrZV4zKx5JiulwC
FtiX91z884aK17qv/jpRCVCuZ25/MoS5ewje7G6DdTLyDW0QXVNNOHtl4zIWt+i1PTFm1KDqr/5w
Gx67h1P53h49AMfR0gxlGITTX51Dnb+o2p2xwbLUYqu+KJbWlK66zB0CUvLqaexOxt3z6pJvebp4
4WLQkXcyf+xBV0DRMPWEiKyCJLjW1x5fF46wocg9vIR0n4TTdALVoFqdgGx/Ixc+2mk3izZnFrqH
JRI64yxVaxYl1v29PscIiv50NedB7MvUNgn9bcXSf+uZmquq6PfwHYRVfFHfHfch993sAr42pgqG
L8o52/M7TQHGqlwagWlHV17ug3h5wtZk24kIIvBrKePHg7uFumq0Yk0Y7h6vT3qJOlw026UbLbKP
IrZDdPGAwTxXF0dt6VF+8VFwNj4e6ZZz7wA+adw8PJbNsF0JSEefC0+agd5kMvIkwe7NitNaLGdD
EPhuud6nP3/+voYkobPdvBcH0oCT1D0WqukHuUgRY4u71nw4B/kDXEmRbDI/UEQRhuCWFj74TZwb
65zMOURdcR0qAKF0m5Ar6/z8NGDqDsgVyHQInmJspTzq/xaFuLC19X2085ZEHTimXZ0LXeX17Iwl
Mw9cWaLVJTcRPPbTVKzdU8i6uoSHdBBl2kCHqNxUgAXrAfbDxluVGEuRWztsL2OEu+xJvzMdub+o
s6rtwHVgRGoA5mRnY5m9qvOh+0u26Vg1Yv8v+jZr9HYPABR/Xxf5RGZfxGH+WbuyEU4N42UzsN0z
nL4ciS1fjNa08i/wLLn40uQStb3GGlqUQblibg48DqZGOEFFaLqQwAP2TpeKmd0eirt+jfUYl3wb
Tn/Bqv5UHCIb7k+/EQXaYKNs2/Milkn5PrSPA13ySPPYxRY+SxzWKrDndFj3DGZdZiD7ilYLqnb3
o100vYemyryFFzivQuaEZ1PwkM0vxk0e7TUKFKx6VkX30eStvfZ/8vQMG4i7Yh6MDJndORw/BtQT
qJVii5DndkHMulJwTNWm0iTY2AZN6+BOb30MpXbHs6rAis1Kdnl+W0zRuKraVpz+RoAybMLE8QL8
HPPWQAR0h08e3BCuWnSCMyP/++DDivNfijI9ydbxHFpKFOdY7f7u9Pe9HsSP6BMfS9gEVbL40E29
9PR3GLzPlCUGhbPLbTKYtPVqtZDchgkd12oULhfIsIXt7zaAcCRfa8yobtAdv1/VzqJyK9241nTv
Bw0+KfqtlHdjbwjURr604k4poJWFomcnYBjhUYWIWwcdJ1me57Br8+b5AOJMobtfm41645sBi/0J
kcg0wkc8KXkyuUiJrR8jAQ2yobaldSu/73E4KafcxJizja60ci8j2OiW51deOM6U3vu0PxilpqFp
Yt1G/ZW1xZ3WvrkB3gIbm+UpkOfYMcAODk94dbm+fJkW58ofnMPFXLXtcsE+TqCRmEirt7Rm70mp
zicWbdbWcEPKuJeGqj2Xa42G8CHhNCX9G4roKI8Z9mALblIpZGuugs+/JpjqcPt5Ocb6EFa9Lau8
8g7n5quZjL5le9VTRaFBcVpnqkH6NwFC2glZ11YgBMNd0tifOVsfsHyBiVnqd1qkQBuEfxFlWrAq
RyKlXbTHPP6nNalJVW12sZmfItcmUdinKhBWxbhmUFF/6EAShtr/d9jPt3qbwcXNutcgNvpnth6i
G09uep/niQB4AQ9p3485YbkPuHk1YGU0XVTLM/WYn89Z3ObxpITsFulu1g/2d0hS8aqwnRpVhsgh
Dfz7JKKddwsbX4eJOp35Q7lrMQYsyn+k1GrAgHjK8t3INkUOa9TBhPpCYtYdvmqMKxWdNfxssxpD
quPkrdTlJUi/s+Bpuz69IzxMrABUfZdG6E/F25+uP8hq6vPK21ctnmTzs/lRcv5rgQWYlvG/3MQz
dTRe0G+eFb+7Dm8tcMniy+PZXtWXeUungKIE+B/Nn0v7RAbVoTSfy6c0kaPC376JR5YJISS0bWmN
95PIWF0cstA6UTGrcu3nV8NHj1BrScJsCh+iYSF8d9VaNo/b1eQLxym67BTp/Y1XstGntlID2atB
4YGvFpmb72UXQlCdeypjuMowBi55O8IFc3+CgKpU15G6VH+Ian1ZJFR2AZFl+Sa1LHQTSiNtCgXk
o1kk0xqSokZZrdNsKOkkP3/sAm+36MlHkJqX/ySRk4L+lRubmxiCMbqwCvD1L++667qJICUZ7/AN
zoqmTIElKzKQ8n8NV3oA2Ldi8L2VbELIbz7QMP5T7fq6SFBHcBocpLwKj63kyNWaeLb+OkNNOsub
EfDeI3rv7xQqZmq6AsakDIgqRe6jtYliWo2KHgDnIJ9OEPl5c3LgBneCXLEGAJwFvLgS4WEX6vaN
18VLH/QJdjDpEF8CVATEa2j+8eQfctc8fmxc/tpAhhuueV17mXZ1Xov2tAIkf61bsz2tbUjsUAkv
LUHnAj8VaRJ9aQ5xTUQDFXQm+jO2sMDvngCcnnaevXZfrO83IZSO9BTmj6ZGxdqJEy3IN1wIpkXn
cGWhP6+A+2NqRlV3ic5xuGlvL3714Olie3rROkhqDpq5tbheoK/KH5lN2SlPnnTADviIg+53FjaP
q8YsYcxuKHbY2dCKHy0ioyFA/55glsNmE32zVu8QCU0uuE2o0DA6wa6AlSe1a8xG32Xo0/Ji3o39
P19K2isjcuVsW/KvVOk3SaM8gk+/kTunAcfpmvwcQvnaGp4sjQzwi7SoBGHsNgTQcqHeQPoIlQBG
mjDciRl4LE7FZ7W5PVp5+j5/P/kWN4DHgzFpWLrAjmoABwxmMTh32qjRy109jx/Wsen6FktJjaQU
1csZH14Kn0yBcM0c/8hUzPCtXS7AQQ506i6ZSrRiwG9vMqSaikXKgrzxjvNQzTfwSwirtl7Wnw3k
RN0rgbSbMmC0jOvjFrWOvG1ReneOEqRtSvmiMkQYD70LZjKfeLHMX0X2J6aEtMxA10CB/x2Lot2g
qJjqIDuxARhPr0t1fjuM5wofE05kmrtf5tNKavSuVHVgqAAnSAt6GD9mB6u2SKUudD1U+fn3kKM+
bWXSQ2adjD9C655kI571FgLREsS+crkx5Lw1LXWTSm5DcyEBLaCMrh3XXon/nyuugFYyHhEUIjGZ
9YyEFtGUCepNQmIZZYOhtmh2/xJAFFVxGy5yXhMsLJb/cBRieTH5o6OybacWv7IXLX7t8mC01sM9
iVSDilvU8gUQ2KHvKbZAP//4gJdM2vTFvWgIYwdgGbjp35jMQuCdyCmrDNIeao/VRdrgCLkP7dio
4VHArY5415gRebJt0ZMx2L21n9yjGhs/pVTWdU7fEFOgmDjt84xUeiavf2nzwNdzEYVG8v/datBm
i2NJIcNGfkcpUdN75etuyNtNyecNfy/RwQ+9oI/NTbqsv/FCxHCMTEyfAKOalq7NmlBakp4D+UDl
T/3ncDE7wVQ0plIN9tfOjkgpmDVWbh4mOXNcRNhTzNUrJb/35XkajPPJXpz8bqMA91sc+uSXhGTs
sAtgbJzNVMr2hWmPlGSozIQo4ZzDEtP4FMNhziD63xNajnYzpBUmQGz5iv8TZLSiAlM1lIJyALBd
r4rcWbCs1DNPKwjo4ke0odOJ3ohXzj3Hroldta+XA720pzoagFtHzCo+1XZPbDFUB5Ie8b+foGv/
UZadW4G5CxG9PLBS/H3JFISI0Whw9532f9xmcLDcrRBjjdet8Rh+THVOb5YfVi6SPsZlVblVOXkZ
TAWycNUVRC0k6pvlFSYLwE1FqoyuYCyrol0BYNTen2mctv7FtP9Q9KI+WNZmFPKvVpcwq3pn3niz
Gl1x+2+Q/+77FOdSgmWZQkLB6ycS2aXQNsIJSN/AhxIPEqWggbb7NQdotgGOQKYLPZA7Vj+YTzfv
AzZzLUbM2Q2eyQv+hJWuNfivASsmIV6ftR+B8nj1QIJoyFv7F2xvnr55PAPlHGqx2thcQIqvqgDB
zbhiQ/NAV0dg4VQ6m3a/PeMVOcDsHkwguHjxV0MYBGPshCX9cN0CtI4HSOtn4Ko8zafnj4P/hJUk
BcEjaIIckmmehgyOCeNUR8uoL+tbMvoK3cgwEI+ysA27NQxhSy2+T6jbWwttNK9EESWrgvxdwa9G
exIkTX2Gnb4l9+ZbjKvyaN3uDpXOBH9ZLEgOy4gFBZnNcZfQwFnKrvKWQPxf+3J6zKfle+Po4E7s
96ZgHuONRtPsWWHN2L4iwVruiQw/jQ70GHiBLcS5npf0NlhRsN5BvAlaOin0EiS5HlZud5t2+MMy
8xZiDclfJS+xWQT/7i2uxSmTfvns4aCRbDPH7m9nT76lHIlH+OWQhKcb8GWp4K+lyUwQHueTJ+J3
WMYrbd6XW4DnwXE6AxVDF0NdHAXpkF0sIjQbHiFDZzqvQC66+ojjZ7nngf+xIRUYFJYL1hiSQe7M
kME4hpfvZRR2xUlzlY+yBh8x/D8wEF9HFnCVdRzhcTPiGGBTHAbAuFEpb60be8ehQDooEXGwS1gt
lmupGvP/KvmgLcelUNmIoU4YpM9XU9lWw98szzAwu/uSAwEekuC09jBxcDcq/LC6GEBBriobnVJT
UYOqu9wIFkI3yQx1yvootC6LJRvgDWjgAHuS7P4Q11QAzNyNLDEOZummEx5nLI8CwjTV4M2YAkSB
sEBgCg/WuV72/zz8v5mM5ggicta4N7JEE0IHqzr8UWjkIiM2GxBVJ2KN7lqtO5t2YvjF9bgrLSH4
pYLxG0t428qK5ESmjwaBWhrCrdgVG6MswJr2GDiBWN3bYaYq4u6uJqmF2y4AvD3iE7qK8qeWJ5Gq
bvENmUUm8kZJhK4LV+jM4Rlj0D5wpfhfqHblRt3nk0FEALVKGQufLMzmVRt6GWXgjSk6+maVW2Zz
rdtBTAxAmEi7kq7aMHrUi3vfhynddSjPT25XkRM/XvEbQLDkYVf1UrBRyWVJgLwx2ZH23wllCDuy
hvbIkuBgcBdGXNrAlpGO4PgpOsEymLVN5IcG2TLYowNXtplVrDQXHeFv2izjCILQKjdID244kuvK
EQNv/Wt8CX8ZEbT9ZgGBiDGz5t1XB0J4P4PNBi1gMIRPe8Ftdc/hRX7B9a76NM9NaIxNHDb3cs7L
0B61wyuci+u7s5gNqoBwFDwjVL4TGKGqAkjPts1ZtyGV9Sl/5Y6diuMJ0754SPCoqMm5eqkF4ujO
iTqYKoxJInjMiZmtDAbdz+RDOeITqtxb5BBH/zCqnq7ebJCrGg9Bj5g7FAiD6OVmyVeKBYjEBIyp
YMlzH55PNv7ke+oMez+F1fkF1Evph39jUNWDvBXtivQFZn27JhfLFcDhMZDveXvMNA7fEQXBm/Y/
nnn44FKOF1DAQiorHsEv33FbwD1FwVWWH9vIcGoE3GFDyhHM6GlJe4OYNMqWy9mpyDOL9sVVt8Vu
Y8Wpt7L+RFOuYE/AUTkPGG+Iy/Y3s8GtBh1Xa0fdQPFzDYXTnZN86mRHOjrBmtyASJXfdB1FRFat
k+HLUbN2inQe5kGDkoEUgJ/JfSHxxYq39ISEvXKpL1XPk3d8orxfmB8qP/sab7G7T2X1k3Fa9o6T
5YV4YEaY7SYTPGfIJuFmCAhGwaVlfH8wwGOEAD+1IYjcJ15LC14kFIq3FKFPQDK1KHWxiKbUvLXl
2H0cZJOXgrj7honhMLJp0m7xehf+rt9YzH8ulxRw9KeFIZmGJidNxJlVPcrHNNGr8QbSRVio+hYd
6YzVjyI3kOhJhxnXznvn10Ir1OB9/KVCuLXHVKQEw1x4yPMwXMsGRb1/TgvCCl43T1tSe3dipH2s
wNEURCT5Q7jULAJUAvKRFSymqAevfxyCQs6mIPYwOIGGR04c2ve5a48YguE6NI9HQyvVEwKp5tQt
Zd+WmLDEI3H83UNvxdc983ED449JxaTwODsLLl8DbDCvaZflq7Inxlq7vIfUx2uzZa7qhdIVQbWV
xFbKXnWs+EOfW5+0zjsXamnyGlemQn8KRVYTE2HXGOMq4KIfsDvVbBeA1D/OR6gH4H0zEEYX5ZfN
47qiuVNdURzkSsbt1kxyZts5VRvRTjaGyVT7B/LOW8Z9F+3nYf+1mwVkBKVvm2J4CcgFppX4P1qc
zShSDllCNS8OLWyYZeVOqtc6nlKyq8MY/IFQrK+9VsZkds/T39sxw27Fj6GlBx+U3kaE2/vreuem
9z0IRtdKASj38QkA3kSdX8J5JNcBl+IFS8mp17Sh9cBmZ07pqXSHmeVG6M+DWMKUFmXolyCLDbO/
uE3CKmw7b7f9ia1+UNtqFT8V2idAPZTxyCanCcVh366beajl5OYWP6jMHsgE5Ac4sWEy0hXqXCrd
g+v5eA/t3jO0EprKqyGF1u5g3n3X8lngIjBkO8nGadREacZZSRhy1e0ZS14P3ESihlNTBQ1wj+gR
nQtAWcM2TwYzDbdNOqTI3DTwqCSbwVhA/kHIL6ADUj44Qw5pwX5El6+lyCkDxYzlZLSmGJua4UOg
8iSAB+qubDWBUqXaRy76F15T/81gPSxgm7xW9Y1B20zvPShvvfE/Xhfa3zR/KkBT0bQzf7uUfOKj
OqoRlEFk3voXmbH5mCrgEGZ5xgnm1lJXyxJ+OwjSlaW3as8f5D1IUparpuVaS2zq7ypZDl0VpDA5
AjSFWaP19VhoArMq117Jyebnp21daAG/Kbxt7SVxOiuwi0INSzGXF3dCrx+uR/qkDdBrNrleV3YN
KkoTyfl2BqwICKYuuJcDk8L21edoeGLY5xwhgKZ80Hj4QG1bNmTw1jyBhTNKK+N2lqI3DCdkj6HF
WWrtYoD5ZXfSzC8vdScGjdp7xiBmGQsDf2r6hda5pUYywtHzRdZQS5xFn4WwvgTTG232EXf2j88o
q3irHoIJSQSe9Z43dbV3j1jFrTmXyCtHz+wT2HLdpDwgkNGmjy97aBp0lGvsCC05Lmp2GnBh8NtK
Yhi/cZel5MLgd/zuyBfJEDz7Gmw8JgAjDCkQZ/bdVK4QDUj3wryjc4FlSBtmhBamuMGF0j3QbhFE
0VWu2cZbmpXJuDFUv1Em7YQzs8RzOlqsY8vrwRXbCiuY+2MDJgCT8521yXMC1k52FH3NSMVlsPYd
4OJu/POhvvHEKckb3WSoMMEuMyJ2e4VdNBX/F5oo5s9CIgvjMeo/paauio2JFVMcq9aSZ6bcz+Go
E5I14KjkgMut/IQQTM7Dpaf37ZRl4Dra76aYh/eAU021NlnUdBtnbDkLi9KBlNSOHa0MElqBHTSg
/ifyixrqHpiOlKwZb+cKEKi61ycZCJGDOMEm55pMVf6la0nfiMzPMRVFmGxlPu1sArtM23SrcSXN
GgDxVDAtVNIcfMeJK0IGoSH7UtRrCOQfUwPa6EXB1UydTsXbkKok38GJwSBH5z17n+7OZfgoQjdo
k3ibh1r3e+j4Yzxom16ILId1aZHO/4qnlwCoRChMtD8XOVpZsGadmBfzS32hQX0+BCfmWAJDV8Ai
9GCKgt7hmVcf4x/R2Jx8LPL58GNfbyzcDOmuhEjdFDGrdP5S5x8P8yM9Sr/hXtm0+UoF7+keiII+
B3AY2XMcfJTIO3ruoAsjtAg5+M6Ps+pLK1Ta9g68RWjcY98oDXndGj+RAKFUZjqCLUUPnn7kTlkU
1qLQR8vZm/fQwHL4srqWvCis0Fb5jm/QeO1ankLUE8U2InXakKYCHoq5N2lSJC46wxsYq0EpRBxC
wQR2hze97HUjvKMpbThplvlxtXNZVt2IjcK6CF9AeeHDeV0tmr/eMzzOt1p2L8TH+ToqNtr285kl
0cuMwpNPDJM/HH3WpoXxKIGoeQOadAUA4usirzJRQdoELFUg4/59EIrSjW+9X4uDOpz1YrWyr1ph
xkrG7jvctaHUE6eDLSkIzPyTJ1MUUQWzr8X8J5Yru7QWwF8KDEwbyRAgqmNf2yQIVpP76QePyYJW
lyNbSCYR+oE1q/DEgfZRAHnWDBqaQE4G4pGvxDSkJ/OMt5lYApHSjzkpGsD13OF/oPOfpwVzS6dZ
7cU6a9Z0G8WSnHlQII7vk13NceKPHanlQTeuNAqGYIMZcmLWXsVWnA2NHdxbP7ofEhRXtM9NK8eH
nublc0Cjem9vO9vQKcqp47tkompeFtj6QdCYgQwzfW4QwlmCV5m4Hv1NNsPzc1p/XwSPLb/H9RP6
zKyubn34gIybC+tJ+Wn2ccTvnnB14OS+QB/DUZ1Upn/0wenNRToY+1rr4eKy1RQ10e69jVfrsp9/
yWmcqYepxcAs1yf6RaG2RJxOSEoQRi+NGQP+opZBmgcFcT5sZenpgMZFAokgLGv74mbvzY/pFe6M
uPlLJKe4PXXFfe0RMxsZVd1bzYcZHmfiJD6Nbr1bNbvPKQGer3XlPu8VR+aZd3pJSzncQlN8TjOS
r4sSLVRSo/ltvJigJNO9MYfjo5c8woRqI19g4NMZf7OGvs75RnLC439JuJ0CGIl4aECTusBXuY2f
rhjnM6py6de6YSiZx1XWptcCjCGv1Dj7EBaJlU4p6EBI/GT1M3qkh0qu9VW/eJWWHrUkztA1+mG5
RkVpr/oKCLMNZpSlVP97Sjb03iGXXTwJZN/TE/Z9UyZR+b+UQo0elWIyBZxK6t3qAKVR7yIaDF7b
++wmNdSef3mAqp5+LRzjwkzIxiVVJ1wzGI117yWDzfkhhJE8rSKVB1IFSgMfsVrjKjNW6xmmIxMv
G8aMNgv1+PS6eVKy27Pkrzfa7BURTbNbI0ywCfWqK4wIn/o6KqyT0XrPe/5gBSZLKCqap4fc3Hn+
1eDp9tCDIEbv1gnpl830e6Ua6nFJmmbDKff34n0Hx/Iyuq8XyOyCPwom8yVbf8pAtfvSv6LYlBMI
AmdFKl/D2pRv1344tomdTB63PdhUP+jbP/zIMqF207XTt8kSPjK/PtLXRP2IHGCHHxJwMPSR9O2j
oMIaria5YxItj7v1snT1VlirH3mTgHOvMUdMVsPVuFUZ2diITeGudS4YdyrnidYqpWZjdKl2t+lm
7LlAohVv18FFTL+mVrPft52k+IH2eW70eDvk1IFinMWeT6parcpbHkFXCPl1iqtQVwciUHp6DbEx
3riY79uQS0wSNgwGOx6cG7EjGPMV/QN0h+7AICsYaRFGj1VR6qfY56204pSouwE6z963bxcBQHjN
o9am0rC2BMCuE+gtxJAb0zGpoSYI/qMLr6Yj8tjTI/ax6LlhcJZoC7rumriFdtJGy+xEc2c7FY7N
l78ST9VdN/dgZMmmVNdXRIQqbDcIcUHMYxyGLEvvkccX4ytjw9jwYw2UjYFu6qAcWhGmAsoWx+8j
FyDc/woVyX9HHEm5nZqHhQSqHkg9yHzuUx+NkmQLRSUhA2/sYR6knHVBlInzfcKC1wtMVEcgHucc
epkmdjg9eyrodlfil8CPTrEkqM+KZTyDtPYVep+WX+BQA1YFClZPri3xhUBAORT8mqqMFNdleOw6
XaLuCyLja4UJOa8uwGAWGsODiP0yndEWtGbRHYhSqFwBfEZ2Y3b64ZxT2HjT+Flb4DV7d5gbadrH
4wsV1gCjkAp5mRHfgSpYO/Y/pS/DrIb342ZuqqKUxClqgP7+GWqiAOD4ZC8Wmn6NXNs+RrDo4HZ2
0pyXPZz/tYv0yow0FbCMmwRzSgfiZKAqDZTADAj36bPok9lkw3Av2S697G6dMcFmBPG8djpirp3L
bESmEYVWqp/c0OXoBuy098JwLkoFnWLrrBdgBZE1m/facw2ATNlfXnPo27vURSGRI3+OFSl/R724
iDnRrxWIlgiNUSFZCx/SxA+ACeqt2M7BeLNqyxWzF+Gg/yE3sWKwtgG976RakIaswsIVzyMH1M5i
WQvQaiCgbDHruZ9Kq63PBTf/MWnIpfymy3h1IwiPS8gYH6hEQh3RN7gDLFOnWkyfnARCP036ASAg
owhZW+PrY7ZCC+xCDgzqShhzomZldwsMQ4rBsfp3YoJM2RWAFXwdZCrpJDvbmJto4GgHB85bwTo8
KG+aHBh6pLIdIrSVdZH1RIsscStWWhG4PoEpYeO5qdqD/mb+IU/FeXtoX2cQZ5QxMu1Kp3UNAQuj
Gqdd4pX9wWXnv+hdJvTQ/C3b3nzFicf1clpJGus6EN+VCYoGJJUh9RUb6LMpZfqvTcfpEmzf3cOP
lHvvbAoBZQ6e/FetjiU2MQkYc55Iaqdt21OnDq7A6QblUDlxF/kV/QuMFX37l28aaFouHWr5DCK2
eJ9oYzqaFQin0eH6rLgfVLDoid7/mtoocLut3BuleOrf9XkZhxLOamnzmlaVPG13++yjbR2xmgt9
lscbrqozT1U4cmedZollIxAIJsYi9doKEUZFTZwEnG8zzi24hWbmMrd6sGT5IOS6dDAWoHR0q70r
UqZPusSCoxqpMHSKRBu5DHxWiTim1UULDBaulLZV/vEq5uZT2nJNmXl7W+rB1G5XPuDkcx85um9K
ED+s0JaPOk2ObSSSsvChYPIDjv6LhPxylJ1I5FIdrWda0kX7rmPXHsw1rrTNWFjtv6tjIU0f5hQx
lSlwh4JqE6Vs+6QCknvR4T33IiFKJx8LeVupl1jjAo3R4oLIQd1pzRBCWmV20V92XKhPHPCKl2Uv
gStenHaTDjBd2e172YfQVSFZd5aXOvlca1q63op0nXPUbgBDUeY6YLcBOPU7VRaczKdMk0K/vG+u
767G+PxMOrngzxOUhNHRCU9bfP8wS/fOgEN+Dcy35PNFqbrnKNh3iUIlPw7hig+JHlLHDZ65JJoE
cOxYa1g3wV8LYPAYQ26OR2AZnSuboIN5GNXLeU4rCBPq5gCip2fKebdpo4MkqFKKnYcHW7mQVvr1
fFgvnb1X4mwTCFwam9aTNmo0qzXjGELeuzEOTNyxaAevENqldgdfFY6FYsljUgJMUvB4Js16W1op
XINcHUn/lAVpPSJFUlbhFR0Vq/Rf80lqkSyQ/WEL1FR+34VCoRxYFazpN1h7BgD2Lv1fFUsF/90a
nvFFwtOjoeybqqyQsde+7qiX7TLJOJ+dpdmXVz7Y0kwRvACZOJh/XftD4YHuIIHferL+KljoZZyP
rwtDvYeHsJcjran47Tcui8yKAofMYsmFZxJ0oKXMRz1g8L+als2eOpVkXPApenJy8PBDJhvLLdnF
zlMFHyOfJjhWZau9j8OUllyJUW8mnPpPMV8UqHHp76SuMl5Ch36pd5BIx8QPHXTw6rJUMRaI5rEV
PGPO8SdCHO8RyaMEzpio3iC7j0/s43cizPNvwDoH0DlY4skRo8pa4xUJzS6GwbPcBbrHOaOHyDeY
X+E+lZx2n56JVFC3a6ZcgxuAH0l11aKm9aUNoIwwuwB1NeQDu6R7A7ak/2FY4dl8cw984lLWxjma
h9mnaGQmWpqwmJGx1GPCtkQVVIXq/WVJMiOrM2RuKqSjhdjD7E7elgAdM6K9I4UAMGRZiVV11n54
iBEYW9qyjTtV/pVholaj0OvDenUguwp06vnOdFg44NkEqXe1LOLlzDJGbuJjdJq/XxXi9igrKSmo
snvjxEMV+5OTsxs4fEFb2HAub9IMnvp9gcTafCUMjfGm7li5YvgNuzYWtDLJjTWgjG0gOC5VuOED
2CPr67lomfSynmx/LZqNAst+iGT3TD/uCgwDsgdp8wTSlGStwXSEhrctD2Mg25CIsMvDzMS9QTsr
1OpjJB8vw9eXEC6Fmgsilbn0fznP7On718JZsQWeUMKcRI264azv42MZeiuUpWddGyaVcS1hXaui
rlXV3EiBLozRs7qZT2IYUYaYnam1RdcHpjyAaKh81643HIikdOLBex8HjLVgLxhmEijb56euD8Yh
2EZDydBDBxs70mQj2xC/DRD8o6FOJahaaz64JP5WPNTw/O5veewV/GwLWfhPizp7L4VTbDG6fNE/
hBgPGPZS7xtMJjWxMpw0wDwH6MRaHwYzQhBU4eeXVle6LmlEO42aBeP7JzBhuiyoTttBTr0ooR9M
qFuckpdc+1A4FXcyZRUiqqDV4ucO8/d1eD39ZUx28De4hRX+qt1OAFo28fScYt+AE3iVg71nWW9D
sGOyJvXaEMjcJDWJ4l0EV/8lwQhvIC9bSgpiBm+rE5eCyyaTNiwIYwnbVV01oudC3d0CCkPLAmWj
i0yiSlTnWI0wYc3Q+oIZn2C7CNhYrK07XtqwwJUyoO86EuGT8BPvZBqRc69znzY1CvDtN61eDza0
KsVviYE1mAtCCdzJMmyRST5VTiDUu3LSKxqOKFND+9s9tJDG1v3tRAQD9xN0GggXOSUsmnIUsCVd
OBt1EHd6CZ8Qyde9jYlpxhDaKGGpx5OOxR+9UabMgYRxesZKqKwVdDmFBSQPP/TgAg4yxUGc65aE
2Tvg1FF27jJymgfh7WPUYLEALJBQaaQdlsQiNCsM0LKq8IT/lfOVxgaoedBlGu39UrbP0rOdbhIa
ptEHUFY3OAYNpv+SFsdOoivpPl6XI0w0rfJ6g0+u/HO/NbhkU1U7sxcbNa9+HXfnTg25EskkPjjH
0FHZBFxQl0TTV1jY3Krmk0kAydY833tUinjN4B4TYviv5iS3zloL0H5JWx/eFzAG0rRDvFABb8dD
5g1pJoaqXjRbI/H96K1xtGtg9QbzCVLq0NnYO+AV0TYOfsozH08YtqWk4/TOburbsnrbig3lqwic
eZmlkJ+gJV29isrkLJBxKxM9J5nH0+739U5e0yY2KUCqqk2mQbU1HZzKzAmD37BHbIKk5DttdbBw
q1l89TaNRdfs+ExLdBGfwR6lZn6pfc0GrQNJrxSIrmU19BEvJaoWQzZi595919lj3iGPVKm0Z63T
4wOertsrWkbsie2pTuEJ+ODqGSk5XILWrzQICj7b+2aoNkp3q0qvi5m1gBB9U86VL8jCCK5u8FZM
ntBy+/fx7+gJnRBz1+d9T2cST3w0psZ5VZ7bMVi1qXNrnUXr2o9x8GBa8aFqwDf+RX3O3E+X9lo8
3vg+H8WFliufJ0enJKyO6hzryevohGzQ5wz+eqYomi7ZVSlxiTRoNFruAtFrmQ04bTHIaEF9vQJP
PLx5Nv977uaoQzfN2zhtJX5Nj7v/GgjLylaFT80UX6WWJgJVPgeTJHwk1TaFoDpmHQPGIYE0A3ir
3zbyHIw635A0x/mnf02fSHuPNliTci9PgigXO8NxGFnTALOeBgNTvhubG2pfYLdibaBoB3s1oQeu
Ml/qbkeT2eqoMcOxV+bRQj9ixmm/mu5f4QzsHsKayiCBilSGGi0c+TjpKQ7tONLU6AUPrcllm6Ft
NQhtfD3OYnqkuKZwLjUH4RWr00ShC5LuC+GUBo5n/WXgSSizwxBO1jHfSMGuqN7SxS0K8oRYh3wW
/YmISW1JzGnql7U9CK/a1WcW5q2CUSiI3JaEmjsr7YMkGJN338QmDlxnqXQ+RA+587DwdtFU535h
5hf5YIeCf6qdp2Nxn2OR71p5dR6sV2QkDasgFBAyCcvEOmeTtJDes8HUKt+zIvIxd3E67Tl7hnM5
GrRsR2/6Cc5xhEqemGvaQPCO+bDudXQZwZh7HFYQcHmTdNh0NdKFWSkEWHWmKb4UnNY5V4PR1k+I
bpPRFpN2BtqGMCSfY/pLMsAlncGBov+CJTXrOc6rUOwxF8Jj2kOTR34AbLz6OHfh9XG5A5Ug+kOA
q2G7R9c44e6zmmgpCWB6h9ajDnqvsxwlV7kVYwxpf5AsAU9X++MK7tYQRTqH5fiwnZJPrDwOGZlJ
ybO+5Op8RtntjYfLaeZnQbW6kPv0zbb7vbqVIBppDzEWOARP8yz8ujj4FQw0BXeGtn3PXNPh7KuA
dvgZZQvTTkICzUWiat20Dh7Z0cVfcbHWHCmPkgjVgKVZYX3jmap+N45/4Z7gWam9/LjFonZq/aNm
RFG4Bklt+TMpK3pa41lgImQ/YSNIVazFBBG7rLstqFQGIYFqRmbn8CRyxBxvmANGCVTLeLvBUhUe
DbOLe5Fa3zZMCJTTGcoN/ywfcW5mTn1YMOv8hCxvEbCb5eDExd3DKIby1QqubApZIoXNjG95+sBU
MWbjYaBkBRzFOAYG0jbLFOi1QqMlrT0Q5Qo64OhFnmZewHbcou4rhUNlOWPBG81xt0HpuWx3jrTx
4V8EbiMesX1Q6Zr6XNqT6wncd06YafOx+Mi3P9zzipLJPXySm+S3rtx+/FaCeeo+WkewJ8UClp5S
IL1gtCPxZdi2HXkzimBSLzSXxT+aK5uf1husaCP6x2u1kgzSIQL27MSZS/VE6FWe90wAvSjx+/Ai
BjC0egE0UUHnQLf6vOMBat8VGeupgRCkKkBZ/3GgYoGmlCIzIpPsrDiPPk7HM3K6sy83APihjXm0
4r4oUhylJP0o0tWyFiOMZYhkhRpcK118pcqZGiWu1oiRPPsVzHCBchkG3JbtkskghcMbf7SdrXnF
c2d1dyhUkRZE3it+t6mR/YyKCdgcqRSIoIbENdbGGDk17t3xR8hxUfgokyGUedB0i7wiITwN5D95
8Axm90KSLa/5LN30SiMX4SfpulhAUpyBj2DYABpp9KPSjI/lZqGaLRSl8qRI2/iFOpdDS8Ayq3QP
sOLWqX8VPsHWv/DExLw0AXjSV8CG8EOPhUXuwJ2crprEeQ8XRwtJPxXSQtsT1eAQznPoXlMIXxwC
03ocZphIAbcr+zNDpyMY69l7K9oWA/09KTZnrUSMTB1YUL97eWUCiUrFPgLPGFbxZ6ul6rTby0Qt
Ks5SPmmOusZ/YrwKkOBHaOJwRonpUeJVs6U8MEFBWkJoLWf5SY6tDDsAI4hLf5E8yQi8PjGCpbfO
VSYIWWxAUlodZkqhm43RtdUXEh2D0sBH9NT8dg8owNx0shzz/r9AdKujpbdys67u83b+CIEiG0S1
T6KZO11+JuBnvDCcsau/JR5ukAnvGvbRW6dMPABWk3BMHo5c3scpwVB/1U4IK6DXJJS1MYBIlXP1
7yKZ+pGZLnElLKUsA4snyZP+gNVgFQ4W0Bk8sr72CAfQFyuJbdqHnJy/Ru361q7ziND+hvdcnyal
ZBpV6Umok/SzCn/Uk35Q0Ev1tP7H6sV6438IrhFZf248LuMkpVr+VcNdPfqBnpNPi3+r4yx6reJr
lGGgrGO6vzCo2k06ELoK+TXD8NTbqa4v7ky1dorfnyMTz92TZPBm3mD3VjGZiOjVLyL5UL1oZxo8
OUPapUXLUjp1oC+Rp+JUIWaRd8MFczKg4WG4zCqGrz91mBa0jOpdyxU/MMqEbLcC3777FxqI1XVa
lrWbp7ITAWDtSzXd44iCuhuqc0uayJwhWrvn1ky3/JYs6gjRNXgzhNOkhLFe9esvXWfqWZ3zutgr
E9fLszR7X0xVwNse7k3+TCwEmMlpk80VRjIRhLpiTt0Dv9Ltbko4PJYN3MQCxiGT7fe/3/jbEExC
dXbxjNIjlCizQDN6biSpSZCCB7howZIk+U7tglMLqGxk+MicmWVKx3ApmRyxBBQQXpOUffFM8Zj2
hTiS1jYfth5NJ5Uh9HowH0N4U0GHyd7dCjOljHUB4xJCEhBTvDN+waBEgEoFLqed8BWnq7RtqqT0
d5hUYMcMBsAv3WyKFF/sc7zt2L7klpKVkrETsBuqa9j5S/MxYWKc2ECZN4NIz0PbRHtJRptH7+8h
7Gr08uM8Kn8isX63b6GP+NlvbGe682M3Vle22E2qbSew3wSHFueJmLJKxuZxZcBiuZ9qgjuK9vwl
OJpBGnKtWNyr0OsB+EP8yJb5c5tXw9p2UrxMyfriPHpAQMm9TWedBtL0wDXSKpQyiZuJbSYLBMPZ
0AGCAFX/w/3zHqLrmR5ZExzQX04GsdsjuSX5AR8q6sxROVYWIpNDts242O99gBSM7YOTBfcFvGTC
WR0Nv4SGvenKZhz/VqQZrcAQHl0tTKbAT9wvup0w0/fCSQ89vTM20StEceiB3Y2bbW/qZaOB4ObA
N4YSOgHnw+M0YnkguBn7IzU/tSpBGd9XTCftiKx/zNuHheL0/sGxuwboUinOEzTN1JSMpiirLpo7
5iceXzzHoRdBHd6SfhnYRov/79c/oG+SUM4U+88BIL2VXMombKM7F/xo+cfSD1IMrsc+XiIpfeN4
RpVgP4DNW+WPUpHb6v5jEYbDDQlhjkH44stP3hMDaoyocAzrqrFcD4bCUmkSC99De53YqXqUVojo
yMXzYWvVvQnYYYcxeAMDX9XDd2lUPdCpOV8vEkskVoNPCWMJYefoXVYclwnyBryJqxMNYSzgVL6O
caUSEqvpSfDtnp+hN5PpLscjwGXyisJ0GAPfCnRD131VfYqJQPR5SBbDn4LsweHaixUtqY4LStyQ
NhAkRUXC0RcaF8nhUzdlGjGh9iTYx2NO7iHtqlZWMlwYcRwhUcnFzfmQMH9vyqIjlMyWrsgQ+RCM
VtL4xA1POUe62sq8v67Il74PCtLJCIL6iN8EkG1rNXiCmBXf0uLkGyCEOjTm2bYpDxcFwMn+iRw+
myx2w82vAkvEEkBnmxThNoDHXzUc/th4Q15/iHKJ5L+nXc8mBCiWzCT0sQrxotZEbaH7MaM9UiRq
vt2dqpRLtYIGUTzK63GRqWdSM6XvVgx1puJWn+/RckoZdKRZD2axtpUceaVKffiSxgwiarQBFu0+
NG/nsIGJweXP7kX4ms6I0FHk54MwiGZYWNRTvDQsKjIQxMWpxz6dMWbCPJPjgFVMdLkFgJHvV49G
c1pXmRGj+Cm/Ur51z0VSX8Ffk5lLqgFfHS8JBoUZHUzJurxBQppxiWO6kS9q7sfpWhXJF8rPDdNZ
tXMn8Qhg6WkCmvlNLK27prAGkhg6Khus7vOidJdBqEkDrYdt2qQw7A3BmBuByQR54gAng3Omz0SQ
Y1jz7jRXaLHRN6hLC6I2X+6Y5BhlDX2PgcBBoyGsZFqh4T1A3As5iBu6CePy/UYOXrPyM5a7Juy4
uqor75vFQUTn4TzfkVahfDqoJcKGztGzLMd3+EQG5WPXoA26VNRrSV+qbwdHhKVyqSIy0PVD0iJD
+3/+dtpzFDYFGakwD59fTafaEcXFa7wi1+wiKNxYn+D0kLJW6IcgGTy96G5DDjy3J8olSDYiuAsr
aWkcNDz7xwEOln2MqOFK1YbEKSn0FdShkA+vC+EjeoAiwKEwBy7zXkIm3aB1oyqrSqdPRl75Neu9
e5vvdMSqM9MCk7k7a1MrY3CS+Mg4GR1Sfp1LrZbcV9ZJi8FurGMclNEuDHWzFpHkiZpTkJAtxIXT
i1qC4YnD0koxNFjUC0AC+K/zmzqMj8Na0IO9UZ1T/RloE91GgCBeKAH04cpEh75Cv71JEdwzv4tq
z/mZwHuONXsR+Oa99J+lRl3JZTPFPUO93ujUM0HF9foH4M2AJIH5uncTPGXOBAiGYyOFpKYes7Ls
LE/tZotMVtEnO/VGda0czsbxWUI7r5Frv3eVLJlPt96ZvvLgPUtG+cGyN9nx65qcEvVlkPB3QnfB
A930DgfX/NnM5Sv1zQ2Vl144boyeKutcAaScdKx2X3rD/+w6wGH1Tc0Uj/9w7kyYXmG8vFgbs0gG
cKAxjON+HNb4GK7m6LHW4HE4rpJBy5XAwastg2dw0weklpb8JjMqZq3tNPrdjyNYXpRViO4aimk8
zbcNJW91u3fYZ5emZG+EAykXMrM1IPmGiw9J7Z6WvrkUbhP5BJihz26l0ixBVTAUO2HupFWsntOA
12Oqhdc9drzFtTUi9NrGvdU/GQtJZyLP8j4Yvs7eW23n84aCpNo7Xp7cgRYMjSJUp2a3aORau/6I
gtVMeJUuuYcjT5P/LbjbQPukTCuo47RoPNn+2AGVIUjyUWguuuulqv/eJR49i97wKEULagS76trD
REyYoFx10lNCkNzCGlRbXebaykdMuCfPJxFp7ERcy7Acg3JFtx/zSE5QuEnV4kFLZaBlUX5xf2+C
+KBARc+8ueiXjgrCyC+qRynR0D6hGNeybxdvxWGG1i1wu/ufL3wxCVMg0DOuCGuvgHX3vn/ovUu+
L2NwxaeFo/vq91X+M080MWMYSp21DFcOcqx+WLk24zz7q1O8H5m8TxVDDJlypsiViqH6+BULHkoz
3Fgzb5HsF+l259CE6fv8ZmVQbmO/+eRkdWHpfK9h6HauBHVF6JXAUT9qRARyLdgBY3OMCAnuMAFz
Ap1GwihQiTL9qDFD3UgFNT+M7W/5n+mgpVIZEJHZTPdODliQ6+gHofCSUStkKea34zDsA8f14Djk
LYQR05qSfx3oCWTmHL8EOB1pTUrQ5Zq01i6pcFJ0mKugu/z+gSPQCDdm80IU4K+58nPDql2Y+Pgn
coaIO++r6FWbYwVcY/H5by7lX14zh/0TJKfLbPsncvmHv+PZoaMTe+zcS5PJDYAK8jdJqDERurIb
iKfA3A3WGev9mIip0+I0ygPgL2HHL6OshdoGwIkfCOTbZ1Z+iRWYofSw4xuLVJD7DI/xeqeLEyAR
+hLL/AC+Uwsv9uSkUhwR9aJTnq+NvslXkc4IvFEAfnaA3HM5YSEXTbfgJN70ri0Q3MDYymCwMyv8
WQ0rD8jq5Ivn3uIwctbQs9Ul/4YWtYEfIQnSvK+w9Kp5gPopAXOEh0rT6TWp2OTrG8J4NZcMDYbI
DvSyrfD8Y6yKSO0ZNT6eDIP2g8I4V9zTO4u+5BLpwXUVQKPUYnIDwkmTMiMXh7/o/WBg2PlTu1hN
Fg0SvPNra/pBWebX/4YsfBdWmQgsk39OeNmQSt6lkf+kr5osxEp0qhb5lgjem7FYA41eRba6tRKH
e1MxhIU/C4f4XfMhy2aKEPCSFSlothpQY1vPfW3x8R10pMiShjDv8eymbEdVesGcdoqGSa98acix
JHL0FzCdMmi/a4SI19Yi5fo3Ynw9/T+7O7hHJ7tls8yU6SmlujlpaCXEsZj8A1Wn47R2lFlo9HzN
oD2MZZgSX03FHeDQrIbJkg14zP9sRi2R5SgvG6HsyM4FtbC9mgZRpzP+gkHL6EgtlYiJ5lhroxtB
1IxvqxD1Mi15FwOwY3MfHxYSC7wouUkMeTC90sG8f9RkHbx6WN+YkHq7gRM8PWg4P58LBoVRiZMn
03GpnJrz7NugBp2J+DOLzTsiAHrX4japJ3yHVjaIiBQBpoMN64ui5Ayi2gzXDY8nnm8C8LYN2dIc
3pym2DFZY+Jl8sqyRlBnAWfgTQcUvVftbeOiWSZJ9Pg7IOsbKvn9xjyAyrce3PRaeYIVCgdAx12W
3sPRR/WnIaH8gEofZsA8bWdC80fd6N9QU4+1WKx1X/LUaEkicWaTrXALSazjmd96EXjQJRqoZ4Tn
JPdzAVh3Z0t8VoY9vYkTzfRqu/N8rdg9lF1vDGKft2fC4g9Diw3K0P40Slq1QIUVpPs0Ju+2uR1n
ZoDTzvusBOzf51GIIM80YYZ6W1CftiG+EGPvbhaPrNv2QvhvNuYYJkotbmqi3T7Cuji8ufvBPk99
mY1QvaRMIGD4JyJHIoEVFS8UfcT3i+Fm5dut0Ys/ot8oels6IF5gPoOuPyTrP0vpqCW0x9I62hz+
zuQkGNTgEAubSNjSGLrkXU027Qj16YWZgMUSokV0jJpP0fcpsDzHEcohG9FF3bNQMNzp46NIzvDy
X0smbuEaR3BESfvaO8A/KNWAqyDOQcK+MEkudMXBPTmdIIXoc3mTYGzfzL/ssRszIxEu7J944Poh
Dsz9z22HrhMZxxMeQWGqtxJVTYQEQCDSemWt6NzxD6ZvV8K/DxcUhWFR8nRBLgmKKTPDdxjGiCt+
h3ccmON8pRKOcNXEy7RGwr7gsDwQnkHDBYaTG8TmCiR7p7w6tgER8S93news7kvIAVKRI4zI/R3/
9yzHOddkfSDP5hsku0sf6G4ga/yT3xwwo8y9uVB49pfc88MX9akzfA65AE2kDIOurJaE6r9TyXvS
NDgOlF48/QYNY1t60EaY1jZb8IrgVxYrPLbxjL3VdHxDiq9wG1lkuN7v+AUmrbniAtKOqzNbHZ3C
pI8EaKziZ7NySfeKNRiFGzjVP6S7D0e47Z7jQ0itAcKOvznI9hlW5km6PUhGOQ14GIic+W/ynq/t
O3RYM+61krlXKsnYuNHWOyR9iPNxr7hfcEt67Sf9Rea0yusZ468s6/UPHTGeVbX/ChOhZvWJPzxt
xwWIcuCrihryyqZ5VJfMdjEoYdUXI00dwmqoIPIDulvKlOvmb5Izy6gVUBRWyhTPjfbbWEL4SjkR
vMeVhZD/GJTPSpsyuSvSphj/NgY8WaPP3G8lEvmu9aydOmoR6GbddywlcMdP7+ujWxZT7tZiT6QV
h51AIyMbSBWzYiMnsGAnGbZpYFQ7L5ZT9UuOHLYRyrxCZ78lCYlhCy/dhlguDm8EtrAWcpwdm8lH
Zmpvc3OcD9+79Wi9yHCuDETo6HgekTRKDwkMu+tre9ZX206JlEX7M67O0J++CjeECI6nddvhWJoz
zX2olGNTKoIo9/fWVa4WyZmviNkhVQuJ22Ra+XLuP06Uhu7rYeEAuNLY0aQDB9J0DBRip4n6mkGo
4kdZZ4wq+EOdXNe4PiBz/i8Strn+Jl9UEsTfsZa+aKpPu/vEU8VBknqKQNFTd7DYzSWYzMpIMBi6
LFFZZc1vn9/GuJ+gVc4Efl8bCISHRaXdzDMen6M9uXgMlYXWyPSuUFhkPJBnWuMdF0G+yVyBA6MU
5MN16zYGBw+MN9BjBMx6/zqwal0P9sTkG+rGJAhTyFf/040pKeBChX+cq9DV9ia5ZvKa1Fhafe9f
yrVR75nC42MnFHhLNmnScqpDS1UHNM8GMa2mU9SHbe7mCG3GHtyr/ZFqCgNr6dUcVcIf7L/XQMiY
x8TTDPE+i+Ad5zTVzNSr3P/Z10Ri4OvIA1OCNzh5wrLyhtvHikV6VBmUZkQoTtvnmMfQcp22c+PQ
jE5suhDSMed//HlVln+JX6LQFGbE35S8JN2j8womtgoX+2OdEmYOwEAPxk4JKS6xuL+YlVKkLBOm
aEMezgm9/jDFPH6Lu2m34K1/+exgBodhGOu3u03UYMyLtGKlmOWytGjLHvkZtsa53askQjJaUqYe
EeEl+oTvmvEI6LY4VQN/p7X7MTUIiroSYRM4nWpZtEsxLcYLQbdkxuWlEWc9bzg6oYJMPyzsSAp4
r/VrtSO8+uLeNpFnrG07PV5yqBTmXar5xWvbSvVrVfXDF1BZOZbJ/U7UoU0943zKvPtQvUL16DVL
YB/9AZA+M5wQLXCkFg9smmFgQglR880XVJ3aNbUpQRLDoQMuAewCRFVP9m0DiYMz4a/NPD0PHQ4E
GUbJ9R7xuG1YdW0x4Q2fbJdd+H2CvvqT4qq2JZd3oonvUuSftcQMuBXAP9TERmC0pfj8hSFmOScb
5KLHX7ry2Gtc6NQPmQZLIoDaKS8uyJgCDmZpJOukH57j4L0k9Tr8XFsjPTCYYrLfSyPU1ANGYxXH
8DhH5e1WDjip/Qy5XUm+hTMrIcWeHdjVgxNbXtZtLJ6PizwU7LeZ0FGR+oY2g3uZEqbWfGRV86Qq
RvLeQEAr2DCkthZ3suvoMazjAMplP9Fg5gXtG8Yh3xd6SWhj7IXRsNC4KK2sgmx0Ov6UZacaHvO/
rK/7sV1sfGNSgFyDknJ0jXwa8b5kanWyzKZmyFoW7hb63JYR/pJfSA8E0OnWsRZ8zJegroBlyHEg
eZ9dZM+5e+x9VCu9xLzYAvo49TkCJr3zp645pjDWGjxjIMAnkTkVxXs0Dhuv9rtCxBCaEdiVXHpd
gBHRVHReknfJq3DK2VA4qYmj/r37u8YVGS25tvU4ANGxg0P6b8nLfJCkqHHurzqh0A5Ub9KPe42h
IqKj1+uDCLXeon33WvhTldD53XTCf1eZphct4QT7YXif5e6q97Yd+f+uwVLTXbFDolloZY12O0yu
3JRcQ00NPdW6QCSFBa3F5fUk7PdAdubxXY8Z6S8dm/l3Do0Q9cNMDr30b3pDxm2XNf8+PSbYP1ju
5I9206QIFgdeG+Zyjr/imNdZqFMQlSpG+r8hCgrvrcdVEPfCATqFjiIg2m6U5uDZeQnF55Ua++hS
kGbvSb8rRsLRuK2RTQAVo5W1oph8A/TKzmChCV6R3KFoUTsK8/Vzr5j/KkBfLH1CsjS0AyL74XSU
ES9bW5UpSZN+rmBQuZ8mihp0UFXXYj4DGw8V6OnYB4ku1L8mTxDQBYwkh77c+rE8K6H5P9nW9BdW
7lL4UdoCNb5tFXHlsZbx7g3lCobvVB7NDbX2uw7As3egln0sLWJotzv2XMjEaHyvvfkpD5U4M5wP
/J1j91Pa4R0XBjlXrfXGSqmCLLT8oDi659nyBt2WcMwrJiyd96AFJ1sjI0n8V+T/MkGBeYj1j8Rp
Dmn4u0PUyXLUuW/FnJCi/fQoESAXGTbA0ngG+hyuKCJMIXK1yfP3DePv/pt544ykKfZvqMIwCPpf
rxf8ieesY5VPiGCQtfcB06KJH3VGJz/MBqz4+/s/i4gJb0tLSnk9gGMMS1WVMHxI+w7FXeo4yG6Q
g7+c6QvKUrgvVYOMCWTMB40uDI439iOfMP2RRd/rlOjP+nP86NYIe0Yw0Tc3amT4p5tZ2FMSApPc
IE68C5Mi6L1D2ymaJIKHgpZi530oUJU3UdQlpiUnQVhUVjLXqB+zaa1RbJ2PoMAwCBS/KEce40Ep
1fJ7JY+eiAiL/EDltV/nFOKwK1CB90KzeY7BpeOk42flyRw4+8rMHCIJ9dcsBE5cY1clg0IFIeoU
Hs4Cq2Jz2sd1r8pVQaXee6ifPI1XrtIPGpL93PJz3fe+d/D5HUBDLLlOZjO2rUi8CLbL28Mlg1XU
Q2Gpujp4F/xMIpF7BOFb/P83hews8vBIJeIhZEEpNeW39OpQ9maYWoo+6GtOfJzLLKomlmknPI0P
y+A1qOaUJWTH/DXpd12z5NfZde5f8twIuajqpS9NAl4l+LLyOPl04fhF5TUHk+V3/ML/c7S1g/r9
QxwSY5eQwTbqgeSx1ZIfZOYgyr/n2KYkn70onlzNqxBv6fJJHDyyEq1AzNvf9VP4JBLESI+p0wcq
6PAYei2yYcxzcsaQRQvc7yaG5AU3jh3xNWX8SCpo+IlIDSSOTZeHeRjxtPd3iGIFGG16KBQlrHde
fKzIt5f7MgpSgN/C6YWX7bs4r946hiZnraNMNoOtpk0e9HCA8wxHQAW999UzFwAuiz5pWaMSI4eV
lmJ5ATbqOhbSjVQ3MVG+2u0McaNlQR6JmR0rrRHRBWGxFPSrCV1QJSwpPHdYHXTVaM1EtQhjWVl3
GwYe0N5IoxXvVCG9gYJ7zqCyE+E1l8bvicIDlnFnQnLhrtihiHAySkKKYtBz28x4JIMor5ZPXUsI
zCtqQDllaRvds4AhR0Ttzi693klCZ9o4pfdPN2khmFZQX4aahw+Y6bmkIdxxp6mqVWwjMfrx/4Fz
kOTx7lbcqcZwARNTqBB/1HcdbUsr6/2XkUZUYQ3Gjg+HZTgwIjkYzkZUAxwT93DXMIJE5BoG+aXa
oatI8hM4wE7XV73LTF7UamJ8xHCfeto0K0Vijpfcdyj0fqB3vRTTxuOjYCweqoFUvlAuTJMs0Ml4
8SzT8xDZAO4FgA37MtE9Jzj5Y5V99d/KM9cLVG+OPImk26IyRRkEzBVxyTjeZxaWS8TnTSXGtKjp
pls6VC+TdkKcGGPTSksmiICPdy+zalVd9dJTFeQImTxUrpUwde4gE3jeKmyR1roK8qCm+oVMQDAS
X7RH3l01zKu19gYLAUVh1FvSy08YAdtNTCBgXdhEfIiiFfKddcLQA1gIoRSjNfrXMbaN1uJC5gTs
8cPaN4QW3szSoT+GFnlDmfEda3Pnm+pozBKyCR/KbD3QGIKS0Wm+gfJEUilGwUEjpqMnzcN/N9FB
sF1RjDXmYd9liEB8F97ICizFzBc7ri6VSE5D9MhjSdQrZGy3BiPqoZrN09hyk7bV0cbjsrjEoajn
P8M1rNIp3IP7hlPA/LRyO/bAnSn2XGuvv60XbCyq1/of6d83W1oIhfAo/e3LnxGDvFfVHgNz04G0
xGUzIQcDdehvX7aSEaoIGBHEjz8ZokLlEEhOajNAWhYAiIyEoLgRj25lbU2MME3crwAuu7wAfSFv
H6f8Yt8wYRuvFvd4BZgvauyWJML+7a4YVqqVMZOkspMH7okg9PQUjDu5CafYHuqIzr2Lvkoq64z5
xV3LpTQVuEM9Hwq61RkBUT4iCAeKweLdVqoAW7pBat914DjluIzFIlkt+Dx2tlMkdsUqG0diBwWH
JvdewtjD4Voj/SAvt86UEJ0ZEGxTOCRla/apgnQOc+uQQily/ZJ3BZEZy4hAMNJGBmIjz5k1URPk
VB9yNEbSKTLYdv+BgCwi/ThcsltkZJtChX97CNhjIJHhlGWP+SG7FiwbustceGMNa6kvOQbVOcm/
OWfH2kcfAdxhJhrgrJvJ2IDX1Jgf8kuFjPPJzHN5c50mvRu5qngnCSV++c2CCBflv/IuxGMD7T9P
jLdHVhxZ8c+Tek8/1m7XGz/MDASy4h+xCR8FHIHCD3cxiYsJmGZn7j4aTi+UYW0NdE263SM3O4lX
SYJohcppQyYeohgUlys55QedlBgEsrxRvNkCq9636cZ7FqFkeuQGhveKQUdbu+lt1vHZnqTVQPD2
7qBHbayD4miLJriD7xEu93I18be+sYmTk8lNBG2aWcf63CXKmV0wrTgtuyYR8exhTUTyob8xCubj
EGwlKuoTwmlEiBqTowJjH4QXZvJ7xDIFkJgaKbZnvJXbpEyyp1z74Ebd7MT0Htu3EswSgNUJxON0
MziXTEodZm5YSWjrqTkA1m2yECNeu6VavAbmOGp/kFfV0FvEacIXsgTskCN9c8T8uNUoB0nIkihI
d0vHNsxx+G3KgJaMVH50HKc+R7ayxfd2K4Zazg4x9iGqZVsa7HvepeVgGJvRCEXS0+vZarLzYoMi
TGa2nWM0LVx0Xsf/FoGEW0m1V7wV+GDZ8qOctLltdMPGc/4Kree6Sl7wr4XqM/m80yf5stHpOsTU
WW5LejCrqIzeIyzMCs5trdsvFR/faTSXLWXTiO63Zs9n/l76Bh8KihlPiQnSExq4Vkj2xkN6Uat8
ULw2B1aZ+IOauR9tGjWQJHNfAYubCaTmKxFuAO0FUhO7lX79z3EMO3sG58CrWvQYVEhIgQBtEgh1
zuoAjStP14+mgWll7RB4zhgws1dRMX3lQs9zPyIQJhsuBa0aptTe6ipY5HQ5FNCLX2kGFMcAGnKa
GW37YWuccWCVEVK1BMGMTPQZov0pXeRx0lLI01PBQH63fUwfUqYQ6kPEcEBbzMnnkYouHFL0FnUS
+ssNKMY+bkPaDvIFiHbwLY1WSHDgDd3VdLjSaeC+U0BTt1DHHfJgWzTJFLkJ9vb2VwHmxGKvDIDA
w8OnU+hBjakA5doxyW93cPW2FkAiNjGx1QL5Z94PHrjet87bOxKxoSb4d9KJmffk2dIV1KqD8xPr
uZgJmFZMOo4Ft/7vg5A9lovoMkZWi7ZeQcRBJjFLqpHSzLlwhi+BVLMLiGl47HF0k3vkcMRC5NCm
R/D6dUa9YiKgVCVMXKgH7TA6k0Mt1HAt7b9uSGQtBm3utLSQd+v0qz+Q6MEzrO12P+tp/zvQkOqZ
1cncUac+/QauZKnBfvTBHOFwxiIKtcr+79Z8D+KqCrUb3xv6mp+IL/q/ThwtfnBL/4MRyQgUAfyX
hT+KSnk9LpRv0X7OM+4YttCC6T/t7K5iQ4CqYRWyp7Cn/k5ydFOSSMX/9yxxw90ZmW2lLRZVNYoZ
BqgjJdP72YlR/rVGblJVU2kK512rp96HdcEqPl2Q+rCKsCmFIgbVovQY1Rb9RfCtZZ+6YD8ao2vC
BYt2oMmOgEmJ1jU54EoXoHYhZ1TBFqjsmea+rOFuvLFWazrEaCeV3spNIaYnfqX2e2i6qzzoLxx+
F7uZhG2KZX1VIjyJdhfAjVOZaCdJc6ex8v6g40PAVxWhZgKSq82Dj+2dt6wl5W8XAIVBE2VjTZj7
H4LsdUD0VLFDm+kWFH2pgx+4smfSuX0RDlZWeXopigE10JVrAVdRtjCv3YGFgbhGRy78DMmM1vkn
crR2z1GJ1EMT0IedvVsnSRWwpTPYgNTee6kR+0FYJWQFSJefzzPgdXC5Hs20Am/dWpeLsR/f07z4
uSId7Y3r/FMZbJrU/K6gtjGSNTwvovDaXvw+a6VCdB3Yn0DpvpN7QB8pHMCXICjgx6n2uCOgWJwh
dWFF9fUSdQKJS/P25lE+M32jQ9wIjVU/3HVJNfnoV2NHds21/cX6T7gN2enaUWal80cQq3q00tct
0j4gDYizQIXMecLhapGGH9W1GsZRfOolna2f6uCVYikWhA6yo6dDxFWYA6ALTfUdTpsJkKOC1D7T
p/xNxy8xbA1BFum8AtwwYfTlXi4L5bYeuoJTI+ezusL+dioYVDbSrDVnYY3iWtuCcuxTAdrdJMg5
bGcq9VR+dZzQ5d+p0eXMGLcPyoevOK6ipvJP1dxxTYTSUyw6jxLYBcZZCYzkWp4ZZR90bVVvDg3y
wnaBcUdAKRO/XBZ8f7bkVSMQsHFmXriNkA30m7ByDtVdgsWL8yBgGl59hu7qFLbIQ/4cuN+LjFx4
rmuOalo1tYh30KFvZ4utMgc56BHRXw1qta4Zbj/5b2h88mco24Rhtb7oliX35N9PEMsniiAyYqGQ
mVRTlu1YnVYp8ZX3FSirNGFfauDYn2T95LMBMupGKh26tNYm8QnnipZnzwGeO26b8W0USjYXFYZA
xuCSOanR9xp3OftsSnAMJR0xx7QXgNtEhivyI0WdCdaIryDh0oC/qXK0/kirCp3S4BXiS4k73U0P
Acy5KGbeYIQ3e+EBfHdZ9LkGErYomS64a3t4+53W5iZs7NVLdctp6eIkJrbbSauk26A7tzoPGm5v
XpFC6+GWRe2muHTlCtuoLzJOkJrt5CfSOR9baOXXnYIA2Lx1X5tJagfi6jo5MlCC1IRwbGM2+rr/
PjD0TJR9/79Qs4DlgCopytmIx1G0LilnEbC9ls+et+riJKzYsM78T6OMYw3An0HYbob39X3qeMh9
Ox+5tfj0GGVP6bV44M7KhGax52HepJ8iBz+Ip7hWWNrW2zU43H+cI/rbzVEnqwar7UHGke7HxG5V
HstMpppAYWNQ6FOzikNkVhOmBaIqF0zNU24u3lhySOnNuNV5JtR3xGuMrVTjgc7+gYtuOpABCmVD
J2qzlCgzui4H98q00lHOrCZvuWVof338viXPrmOFiLJIiTlfTthTdRkKvJD2u7e+wjv+dYLPe2p3
hoPGt5psb9USxOgIfD4pPXUZJMPeNrYV9Ziv8ibUQPJtX505xKuMCHzStj2Enft29x7oj8EUOejO
BF2hn13R+qdF9qtDlvtUEYQbqzoog7R0sJp2+A3vUG4S+aFRI8lLKS3nj5C6EH1kA11adsjD365w
gfWaTNQGKjpSIucxv3n8ms4LrvBLIm2kXLUDemBeLBoDdKA5RjBmOdRL3K6ZgPGBiFg3lL8xl3wT
L/nwTP62NkoPts7STkFsPJRvVbpPKsTsz4ELb7wY1DD12oLTiVjQmyGK390s1KamwQtblhtQ59o/
cMWQSrWVh0XM9JSRPgczh5/CQOCdxH4aNu5W0ftXrvHjSivHHGsEtq667oloxVZiLa0myWkC3OUb
WuDLAsW/I737JIuJ6i0FOJJ0nkYzd6FFp5ct5ZU/qqFddbbUmlQzrjpogRSpuexJmQn4UpJku2/G
ieuV6u0Rvew/Hed46iKAuoHoUYLw+p58kFxXAb5002kzkzVW3zu5vy4bqy0q8YlH2lxWB1uoZgUQ
NamBp1w9Tai3A8x0Noq9tH7NZh71u1QeOZlB7Y0kAobY38IvvGIDo3JTPcqrLyalAA7AdE+vgs7q
TcETOz3T5VbGY+A3nCOf2vqk7WBm83VqNOMJRGfAzDZTkD1oxmAAyDKLR7GmajnCuLnPqBPoMD7W
mOCjWfzpzl2qo5wkhutXobTQJdUJTvSYcxN0N/o97zXWEpQoULQa0Zwwr858Beuf1p48AYNUlDeT
BnYuG5WSexmLzlc96TP94z0p/thXNfk6Nxb1krpNpPTEkb3nqRk4OGoDH1fE0lYvjc080pWGBKde
KWa5UcSWEEHQHB7loYUXFlXIU5P4uo+G8NqgLZRgfD0hVSHRj0Y0R6ur9eRtDZnegt0QpI4nx38R
V5TQaciFO/TFLlCB0pdJvart7tl7dLbYilmsAIsyrN93bY/YbO8t0uVxKhMHkKsExkzkbhah/U6f
hxseDB7IqfVn/RGyOeuRuEp2/iQ8nqgZ3f8qYYtdbjoYe8mUo2mlCgfmH626D9hkIRXHgTsxZj+o
iAV5e1ufxvq0ujAUTaSey77mj14lLXjo99fCd5csaiZQdarsiU+zn/RM9tB4S8gNey7MwsN3TFdU
x4tuQLLSfB5iv668Ph/H/yADGbDOu+UkknEynEWo6HB6Nu1Ozgzd/0Gf5I88ExwEXY1vhTmG6Xi8
cmAHfSYWPbmb9o8pnCfo6WiKMnwE9JY+dzRiSB1y8SpWTdTLIIWloibb3kFGaOo4rHe52qARZ5x0
whvqYsz3QbJ0Nm4bzdWSubEzqyM6BBBFqdm65YT9BycMvhv3jLLlpyJYYvJ9exeBppEOJWonKjd0
tDxsAKepXwFQ2fLHoISewJS85V7EdoV6QQWGZHOqGruZgBh2WLKe8eZa3l1jvmpiRtKHWap9Gks2
vPRsKXndxYeA4j5kvNBsmMpq2PpzVbrIhGt7qYiGMfQfFYqGI10FtwdAe0lH/UunsiSwWWPQh0T3
iEZ4nb8J8bQb8xa9sLwq3+Bekh5o17hg7go2bkZ3ApbgwNRDg39YxM7U2GRkI2iNGWNBFxvqhFOF
8bs489GGQDiT/Qq9cF4Vi5PiJYOatp1LkhWB2E+J55Yy1tBNPvndr8ypxp43K8WQZNTSx9e/HdXs
cQMpVtTHaFLqARkalqJrkQS0v6sOmCRThDk2NBQuG82qPWMsGwgAAItKy+2iy+0t+fJdLx4rB0S2
u52dYZrRXCXSxbIzNOKIAoZXyPHAmf/JKvh2I2+HtJzYXtDz500GQY7TgDwtm1TbsZdEjbmPA6Tg
mQ1aCrgFcDjaYRCvrbdIQivbOMtBwHweCFX3sf7+9G94zuDN9j23Vr3A/2aZTLXmqzqbiadX0K+q
HspCo06/MHCLwXM1w+S0OUzzxkHl3qnW+1TfNaReHkYr3aRUKU+BoOIGNzIOsb1Sefysml4nqo73
Lsju8cS8sUEkWSo/LtC2JfoyZEAMj7XVK5CpgJdZWDHyTEA1gewd3xxAaDL99T+Sdmb/M38+7Moq
dpohTB+7eYKGw6n23QCTFZqqiy/SBz4ZWF3UuljrpD86lhypIaMdnxHX/xF9RT0k04x/T1GBUlia
98BEdsQNxI5TwWzsJLFEGnHeTxrefMMP+M/xiJYgASj33f3gpsfI6rLPK+RzmVgckGr4+fU6wnti
dLLE60kCNfYONXqsspJeujJ85kMq7rxeNfZeChPYDFZN34L2+/snzLD9ojvDdZh11l0G73jqNZil
v6XeEwLjZTm98sP14wdjA/mJqcgI3v7kn4KYqjoFp6xq35xPvvkK/sxaF1oDRov8Y9Ms9be7Qk6v
fz49axZ+70X901NmzzUHtjmz6uQDzNI616SMLfQGLGJqEQeU9FSV5BGiueLviMj2b0CEGiPbG7Pd
5bm2vuHZBDzxeSricSMZhE2HQ//D7AkwwzvUFFwa6GAtLN1ddJn7h6cu5mlSrTUdmfoXWq24mNnB
ECzXAziwVFnA+PRXL3pZAbPvAhxzTgvLsiDeNDHwykJbNmwipx1FOXrxkdfaMQc+8W9th3ZhTdyX
E0R3RW2/ZfHORIVtA36GTsQCg6f6AV3KoCMAxWqAJD9MM+d4B7+2GhQuIQKpLkDW2oHHGN/oMwhn
XBpDbJYEJced6mpZfAEJbBkAbJhH9EGRsZsTn/niPACfbasSOhpCpipDbPs1OMarGv5ptK6SzND4
LZN/G9bkKgpo/4mKLeEClAnASr91fxc/Q+XyCxL/PNPo7rpSoxFYuEtI6rm97aMjWRj04vpJCXs9
zENmWmCAd43mNSAbnOVL76K9vsvx7i8MCgI7AxeeR+xyMGWwBhgAYIztZzWF4X5UNKJbanIBqt2r
FHtt3AEbpYQnHea2WWVAt/Jv4hKAjhoywADyKZG7MEh0HOvLXkuXH6veoOH5uwJLK1ob+VYH/VJ6
DVTsBC6sBiM1CIwiMxFN3czwuUnyPTMvLQ6iK0gGNiiVan8NhrAe+7UjtYjHlX+pLYM28EDthlGU
yAF+vAqgmOOnykYavLXjmFWO6hkFjPws4IpK+HhY0Kyj9cr2oB1nEi7Cr6TIpLPuKAnBQ2XKXGgc
JB1vONCuuJN+i5gRC4/XAszw7WoP6NnvpzJjz3FedDIDiQbS1ThhE+ZWoUCPQIx5A5LpxaqKByEM
SL9vJQ9nb4O3wmF7VFbqBlccO510xxwKe+JBmzsa04g/46RLIZjZQyPt4hA67ne7+hmZCIMLA+ic
TCGHiP7r6FdBwOjmwL+y2/S1uPllJzEXtQdXjendwCh7OLFjjusgDqhc4svtFVTG3TcC9p02tmNH
zT68zXsSymjzJTMqxc0L53bvsMu8H58nxYR3ddm4by+Snst4wP+2npM0YM00ScitDzalFW8pEwZm
9yvJC4VaHSgM/PzMmk2k+6au4cJym8GWWkfL1gYKU15kTnGHki0wD/xFsfHy63UQDaROiUCek4tw
e727Kkwlf+XZj9B32ZEmymnRi7Uum8uKOQAdNh6Z255yRF89bQRkGjulfC5EKqKGZDohlFYT8BZO
ovXUofTmY6lWUYAMy/AJv3MCfMy5WpdFl15QyRNG4M8Q+0rAgEy5AKPh4TOu9VNxr+B0eGtG2M+1
f3NqD7uZ9V8gnukBAlybJq26PT+xPIQ77VLdQcyh6V5QpowBzpPgxJcH1HG4ECzCrQ8wChwTNh55
L4sIdBSEyMW/kfukkBH0pVVyb7SaL4FJBy8fELU7FN2M7o5Y0jI1Ik6kSupFb/q7OGcTJvU2qQr9
V9xwSjCF4+85jBfYpeAOWHHiGBF51DDboyRq/yjHN+cNJiYDw+YukcyUIpsKVwu6n98wuWWcSzLT
lEvAwnd7gr0yld9xey/ssD7edMmRlxeH4vn8+pgfFQdUM+sF3uxmZimaj8OjadFNoKA6g3s4UuSH
C4hG/q37xypjpe1xKRN+MCmj0ZMfLLZGT7JNm98E3lX7GB1kk3iOvJ3NGpvhDWIt6cgdr4z16+4j
+9td3s9MI40v4GMKOvAdo4MTWx4NCKDPkfGxJdD3g6xd3RbZvHVT4enB5ncj+LyJQ1sVG5nOB7B5
jOYPXwlE9I9OLh78CUsx/RJFuXzft5Vi/y5fboMzsGK2QDwqFatw8jesXDgkKzXDW87ElPxmJzNb
L4+HCylg7RuxCUuDgQDkgLXzcdtIHE70VCoYWzjobErk1b1D79vcv6VDpjvvoYNEq1xB8uvIbBHP
INWpVShVe1LZ32xye5qEP2ZHiXRZtXUtFQHkC6USGO/BqfZa9p6jkeEnV0sbFpUTqK4QhJGlHlYu
RH1PhipF+K86ImtLfsTak2jkLdia6nNK//iuefuB+6D3orExUZtejk3J0kEtc2A+0ew1L07VG/KB
P/lKpUghpJwKse+gvjzcZbxgiHDj1f6ZhqkG9p2Y6Nxdgj6tcrUhnT4zOvELE7ElzxAN3Dp12708
82BpVyvlzqbwMJ0Rhn56kMU5/rDY9PxjRM2fCz8jAeoD3zEPt0i4CPARMuyBdcNya1IBNaQWyW+a
TYSnJjukTHkgVPF+aG/8dJ7HgeIq2iKfgpvw1e6TQcrK23aKONCBej8dCeY4T1GAg7ZCgBYxWxKk
Fqgv/qBltrdPrW9v4HUiFRpL8OR4fZiYUy8NxKi4nvqysn81s/ifLw9S/IkyV4AW6DE9FfbsTbVe
/Nnca07ynWZGbUM9Eyx4cvz1nAiVBdjDZd0BH4yqvJkW2iKYjP+nz+7ytsoD/UfAl08jWrgfxPaS
oPDIAJA3Syy7I4NGHIKUx65dy8ZIE3Hv4mWetPByjzG1US2XIpDRREfMJw/jiagxRA9yZQ6wgdgr
M0MA88xta21Qe2S5yxr7ak1enVynx0VxjC83jv9o/34Uu1vbiNH0BmxPgSXe83vQEBSdcYr15E3x
4/Gi70duOjSu/ZA7w4evqJ0MEbx6XsmBscnUylBkBUt1pFC8mHPbiJkjC9mlvO5dwEduMa953OyS
AxUwx01+k2Ivuy5SJZIBYyXRA8dkP1dKlsfciF8vzYQ2gdjxahInB2GOKZeUI7/2QDUyUWycFH5Z
sJ7dFEfwiMz2HfS3XxQZWh3ioO8X9vLuYRFIfGIZqMHSbKgMqok5HDTD+DWkEof4GCWosP+P1Dtc
yH4Dsl/VNvhlhGHjK/RxdR58L9XIZBh6Intu4L+/uG7BatLlpxix431/dDRgi6neM6gP9U4H0aoG
+ihJ2SrnvrOZTap7jAwcBt6RrejMWScOB7FOeygywZWnp8P/NQ901l0HKPAUPTk2dBBhHrQChAb0
817YnGozIszu/wvD72UVuFj7zJ/L1F4HmjP3l3tNXJDerEXolG//6BYSpNXV5SycrQ/QcLWNo6M2
qjYDN8qG8TzxPW6+Fp/8fk+/pN9lvpNAKl3C3DkI/7DLWX7nYIgUtdXNFHPJLLO6C30mee7JZeat
IBSsNW7M6sQRgmOofcev6t/ddYwsBN7/NF277FR/b2rZ/e8EcyGbVmVyC84/WsdRXOD/yn1Teqhm
7TqYhD8YWW3O1+axm8nI0gaUKRteadz8FSWy0THolJAEHENM6jzCZhVq6Tv4et3jyv7LT0TrRPAv
Hlhc2SZ105iZEbrRA7FRyvbQGrr7tlrav8346pOaSsdojPtFGrwyPqlfeKceLEnBCSXCGevdVMFY
W5GSDdimBObaRQoqm5ipw/rgyiHCTYrikVIo0FjYiK3bsp98SWnUauezjs2us7CCepmtbTkyEIdb
goZh6r8ml+WVHPo91k5t81cfB0NiFr3Mz+yW2d2y9anrZNJFihdEZJZbowmHZEZtDEBMRw6VF6bC
DqjSTEtQ5ZJxSfG+RoPyiISXt+80TIb+2OtY36pGEeUz2DsTYQXEm/2t2FwxRmGTC3cF4sck8KJD
T18AZdlOedjFROpzxLMbPikmAOps6+7T1X4wOuv6/aumXKwFLgRubduKSW8j+pvNSmJkZQWYyaFu
F8Yt8PTfy9oWsQ5oMK9MOZxgCn5gX9K+RJ5v9l0yPF9ANmMKIQP/dD8f/CJBzrnwx93Uea46YJTt
WuFAEn+sm/ZWl6cd9D3eNOTxFNBtrBE+F0GC3/iUqWDcwneNYTUkuLWC38PpQHpsg6JrfFCD/6yv
pWkz9eMIhoAJwZ4FS6KFKqFiTSNXGgVZW54JsGTRqJ6WiXWMNzvf0D7vC6NrolnrFr46HU1i3QPp
GgFDzelxi+wqvBfhmNWwJIC1DJzSDa1ua+9zBfp9NA2XgeaTJdA4FoKqAY4aRsqwQfxRt7mlqyit
olkEv35rFJ4XSHk3f6sYPoiWcg0H+ZVjk2fAiKz5OIuhnZH1h2hOQqJSe5ZeupEHXFqXLfepTLQZ
gJ/jmk2JVfd6gw/7bIqRnaAhl+eVmrfKqjK1CxN9Vl/fvlOuBQLKfb0+9M+C6hFJ/T22Bzb3M61G
gmfCK3/R/hl68yAI3VHIMK9tX3iEKMme8tWX/Gv82GM3iIQvUUZOnxxE5K1U41VEECzmEqPtiRN+
zV1YaPVd3cm9pqpAgwn6NoGrD33iMqQkQHL8bJ4fWLkhdPeOiLKeQJqG5gjamvKU+NSXcZdWTd3i
UrL7ScK28FLWztkjdNn3UTMXz4a7SOppmw38AfszXJ/+cGVs0voekMT6O5gIV2kjQxcmN80/T2vP
DkRI041Hai3O6844oZ0PlyRT+8EuHWb+tinisw9gQihxYE+nlSEYu80aw7k9Sy2QFkdiV2nd/xN6
WaHsWVpuRNqUTZCCDRfvGYPriHqnyLByvyzGFHMoyROz3+1h4SrfHcZknCuB3KOJBbvX30FC6dCO
l4hWmkukbRc42yAga3PftJofpk0M+Kc5sdFfNoKeu8hFtjGBiDFHzM9PSe0CFtAnCLF1LE6D+9vT
Evb5bssyyhzA4FBtUgd0hwiD5oIoUz4ZQSaljhrWoaJ+wvYyxE9KV8b7OLRO9kSkMJD9mOjJ4OTV
Vk3sT2zOSe+8gyDihAW34iHrtVsg/Hi8q1xKCJOVEgUXmr689kg08r9Htb9szJusQToFNwTztGBd
FqUyj2bZZNBakI5KfoYLdXbKKrtkKATDi8ongEJYErSCZeWJej3u/mGfV+eODFz/8AkzGA+CU7bu
pAXsNDrjYE6DV61HSrSqKs/f3l2FJulkcmkkVWYs4bU94EN7YIbo2B4geaMzmA7O80+s5VDBeY6E
VBOwwxdDJl9QR3//jn6QzEyfrBN5ShkfsQBDBT0oAbWj1UTZHocoV6A7Xa7Gt8mjmvXBCJ215QWb
HyZz6Ux+7vpScK375s0TfoaY1KdphDETX/6l15q4cGy10wBzwdp8CPQxtGmqwOntQffS099vT6f6
lIuMx7/D7y2AnHO1ywy51vPUOwPlVrFJ2mcQntZd25LFkyapBTyCOFhcXOEvbFMK7DQYBIBjPoF6
YXP7fK+pAGzTIbIk8ETk5ZjnUJtyugqINACozScvTL0D8pdxeQ5KaKNwponJeUIxQY+g2zSCEpH4
vHYsW+Fx0sbw0SDBXRcrSSLvaVoF1EiE9wG72sQFZQwvz3xWTqFGQcb55XpF4050r5dg7b9ccJ24
AUGc6CJYKNE+qUr/wKzXPQospZvphvjoC4J0Jvm9cLmPnH6cIxC3gBg7FMj6Hg2KrjKAdRsgST6t
C7XlVvJ2sxsx0wCqMrGmX2XxlTUe55PTUiL89+oZNEJwZJ3Vx/dz9cpIUxGOGWV0CGzJY9nI/+RJ
yRhn1H9lYM6KeYJhtDm/i55vLyYU/kYhrCE5EbpgkgHLOx9AgYVO63QWUbgzyfqE9QFsFue1o3fJ
eFU1RmADmw3cmsJ9K4ctPT3h4JKe9N1IpDWl6565FtTbTrnOdxsEFhnKF6ceHV9lqonm5nXOYjvB
ivebPebj2mnmAtdH9NKQiDC2rZcHciaSm7f5gXwUXCVVan++PwtenRCnur5JJPdxMn9CezFkN/QU
OLR7GhiI48GWblr6wb9qoyN1a/e3Z+PCQup4QpiYSd2I+o5Wrcouwhyn64sMMciBenXb3eEc7tms
EHllkiNCbUnzwbHlEgcv7zsjgDH4aLhOMolR48EOqp1DwHjNhJaN4CBT6lF82f3KLe5iBqrB06Gk
bZzisaMj6WVWrAbrD9DyDPv9b28pi210nd+NPSkP12aVcft0fI22cE6vJxruTP06ZNvvmbcU5BWW
RZ9giLTO0NHzYKPdm9H6P/ytl9HfCuIIWJOkMWd11RNNY7mIwjRwo0/OT592zvfU9q7YUBoEWD1p
y2Mn5Hi3wg6NVnlhjcL/jrhSn4zv5MM+KUM1y/vfFc+2R2SypLqiLuxxxfGdCGb59rcMNU90Oqzc
E18LdhEp8YG4fVMGPs2eK0FW+IssluRSajawyo1SRLLsK8uP+ObtzixY5CnkXNutiNvuylXM5XQ5
OSgNlbXxUtuVIjHRDQRTQmtSKI7xqOQj2ArxUiEnxT3g7b6/vEznmS1OBrxvzbqUVZS7YzMqOLEq
0Md35STtNm7Fj/mEfBS9Yx4HZZBpvVn0HyxsaP30s20Srw7xzaEzAgMGEl17ymF5LY3zJR7U3IlJ
FhybdnQ9ndeFj8cP0ICkzjjSlvuopXUrpCHGa1sFuGNFilR7rsVY7wHl7AFU/sv2xcmz4wPyV/Is
Do0p2NWtm1r2vbP+9p/cnrsp+obK5cwEOgz8gsQjvjcvQX5fqP7v5g69Jdlbsgk0vsCnSQmGYmhp
psk67RlplgXUj+ZO9FURQIF3GWQHjNp2/L4LywVaLXaKlANdtBVaf/uOpxKBFOSoUcRYysXi0zKZ
VHE1snWQoNv/82NU18mr7SuLp1RI6Ltp2X3/oeUZDzjTeV+6ryKlspowk8Z3ILrUov7Pmb41ZWgf
ixTJ5a/8+EEbGdIBSMHSm1GqaX+TZXTzyxZg0HQjNgd0m2kA78znY6BThX/CNzxQuIhpGsAfdAbG
TlXJl9vMItnjB89WtmyQnDWmK5ws0LByUVQTvkIhcKaNXTaSngS+CSUkL2+fTzzqdsitQlJREm/v
czeChjELGL5PtoU8ZhdjA+CXYNJyP+J23BuvY2tMe5iczOUB3VtDSf3NXkXqLmvC2UfSJjHVOUZx
zIGp5z2z2SmBpbuRYZqHbeUma+aA87lhBKCmuAo8bLrJP91ddfgsFm0WrHo/+L0083TvptwoBAg/
4IITiDoBtXE0dYhJ+TwY6uVQ0kBCXaGeXBJ4cNqIqmoAk/DTMaTcpn5c4NhzI+xtdlxuvCumlHNs
JQ/1MNf4GzVyEpgX1WgZlI67FG+6KOrkIHpLr0raQUTSFm3xkqV8f0Lz+DOPABbaCy/Q1nc6Mv7T
Uwz7kJfrcenai0d7EhPvkn/f0trgu4k0bLbypwZaB+JQUReKHju5mYZ+kT8g66kSSH5qcKyth1Cc
pNgS57uSrkJ2sCawnwanBSGRifH6D6fl+Y6yyKQXJq7IXyTubc4gEsfbq2ZBfA+o4SzHAFTHqy+D
C3GW43p38erccSrtnDNWVf0fsqZwIgNmHDSyw3crCJdaPC+uuVcJwoeC+of6s4IjbUnhYsglI9eS
dBFoqUcVUM7GPJ8OV1fBDFzPUZydCTB8SCnoWMSOZO+PH3x1RD/eKkw2EwqvRcKGz35L2Te/fkvA
nAFtG4Gik+4IYHA809OOaQxWA/1ZIvqcM4Erz3DRbCPXTikdaI6clUFki2Fn3KssgG9tw0OKGlGp
diB4Ot8ZIDMbnAdhSRRuU5NIX+n/p90LuIE58F/oLA+WlCtoqXVzXI626BIZb0r2VwAvLHD9kew+
r83OBySeDecLnwY0HAxSlA9Pq3vw9oYVS9K9Not7Olf7xQ+oyLgdOqDCAfp2zCQCDLOpw0RTnp0Y
ZJHcH1irSJ87jZeZD5pNTV6HUSRqUkX3HhbzLpnbn5gPrH9jsf/oAuKhLEjYJnZKm7G4CO0fTgua
aEAaruWciK+J370qvd16hbhriYU35232hBRPT1xe0xtXduYE9TUk6rJNHTBG2D0b7D6u/F4/wDyB
g1JJSfqiZL57GOeg9m+6Dm/gzzLEXDXvOYkfVmSELybefepGdiqkmqIzcG0pI++rdb992qJgxyoD
bvXWiJaLE6nmGlJDAmJ3HxHxUuQU4z0ccnWWFCPsyc1kG67RcDeoc2JZYQqhUWzrYVxLxepaCMLZ
mb8BJz8xiUYNVRrgVXVe3KaxWvq1t4iePjmef/6PeI7DJ+ldqIXmWQDdE5M/BSIZdlUz8eyX92R6
epBGw04JeQv2YSEtiwEYcCTFZTiby5WwSF/OY+RyZyISkgVgMb684RjnvlU+D9DAJIfpnAQR6r+K
lRK6yVG2yqT7XJngI5eNcAO7KJSbbVeh5dJGY3oysAqu5QB1QohZkQQqu8CpUg8chedrgXdgup6y
XZ/blcnR8lXGbAqD926wOjx2YPjFyp/WZojPIXe2ig0rZHbmJtp7qfUHLFFQeYF6CprKqNobxqBP
tiVK3HM0twex0IPmGg5nc1lDDR/k572PzKbkCJMrU4/2KC3lnaedEIsr99eVZAWAdvHnrGMiG9Qr
u+GZMZpQzzorCig+EcEmtPksNdb7dkNDpNp73Tz6DxvVdl8NE6a2x/VCbiKXcLrLf2V8OuEXWYOb
ls/8+8UiXIKpCMPxRFXzIzFNp93GqhLifLQJA0/+Mj3VGahec9MgV/WFL4va+RMYK0x56lTZh6mN
hedV0eNaqIaRQm4x53duuIQwW/9zB8zDuTzStiJQ58nMLJmxC035pqlUGuwBEdbohg7Y2lcqNFi6
LEkQcEgaE1jpRcatVsc3SpcD/6VKD8q2rhq1JGYi5QU8v7qMQ5JFH59MlJK5r57IuTkcOe7NjrET
xWB4F9wBlhplaEfxI8x1iJ1bLPA1foS6SKyUfRnCieFL3UU1LtYeKmLyosI7yDUGtX8vdeuWiQ4Y
b6PxgNls25bgbbKn6oTkFlC86Itif6DzuOv/fSLtNW0IaNjrqqjDhj0JWi9g/pj0/RYTs3++r+KD
cuk7PvfeC2q4XqeXW/+61F5puAaN3jRwqwIPG0Rgm2NvmcxKM6zXsjmnXdf4RvCT8gXlrrdKMa/2
gsp8dk0kw+MAphDY+olfPlyQ/21n1xLSw+jF8oxdaRI/Um6YHt9rQkDoR8/8QP4Gvhjs6FYtstOh
0y5TQs5b2dK/KBg/llylNVvsKBDJtXtUB2juC8h2dIL/abnooEHAoU728IM+HzjWEMSr4Xm3NpI8
MWzga1OiJzEedFBPXJFYfrmGsoW0kvvNvQ23jOAY5glxTvyQri/6feoEvu4mhTllJIIggHvToC9m
8EplTuUtYzhji4Hu1jRytPD7U41hUxEnd83KKtimsVkiX3XaJ4rGrLDiP4lIzCMYX6OwO9FGHceP
YlM0qdlJbSsZ75RGxZafQ7jtqyxiWzjdayWJqeL+92Ej9jWBsojaJcePZYOW21omTj2NxhPn7FwK
0X+EXEDy105DcAf5pE5i+ejCoN2SCSm6b4C4HDhm+o+zb8FeJ9jLrKWHrMmk07e4IikDd+7bmNol
hVSVNwq/BJL4midC17BohunbVpQoyTuCMrBAkSww03H77Ir2LZbpNRf2yCYXZpVAAwvq3ST1CSzV
kqIZUYxFqk07E4SjIeTl+2MXmGd0MeFZYFx4cSdnKMEXDmlKavhzxcTC61nGI4/aCkjw6gzdfid3
UNyIuRDW+K3lJj3gG1NVuyUT/pF0Fzf0HzKWAhZ185SkZBvC259i/XwRH0Nu1ImEox+theyqBSIW
ybOKKc258UxtB8B8WLVa8tY7F1zft+8yeaJOjoJWarYWsi8ehaw9atOvA4paCm9Ddzaaw5BESOuX
3DE+Bs3o09S8rqCoz3NreNakm16wMCkw7PSXXarzbNUIzJBspaycsDoDkaSVMDVmBHuJ+hQkIGoz
tOargi0WK8o5ANCujVP1ZJgoacVfvux4nLfylA+ixMCgtjoM3RU5H3WFdVaoME7/mr6viRaCJDJf
vp/putLUfKtLcDH8//j54vmWqiG1tXmcsuk9cM8/9+s/PrvQMKLVPsBMo0BdFfx02N3NKfZf0CEz
K3ln3YYBQ6wfU2VaBnMCC+OnuhlJWqMXG11h9HCjSo4+F3Yo6lSVP2SI7JYNi8eg0XM5GR3hMkb1
jy0uvYY9anQMKEtRJNxA/RWeixSBAp/q0nKf1e4JT2GmX1JekCw8uDW/ByVSoVfcBCpJ4Fb+Db2N
FUL9cCiI1W2bVYzZ1Fw+QEKfU36a9X97+J3JEX7IXanfMwkdW2Mcn+WdCJGoy0MyK6RiaFK9mVCm
8IKKApF37H6g4ZP5tUTFUcH2lUEfeUG4XYd/dqEF3ZmSWJeBSO+IL71jlWyDrqLNBYyjDfDkcbeM
HPcmlagDYf6ANHBfxO4nvp0/+Hg8cmSUas1wPljrgRq3FyT5I7JbeycAmOGhBnUP7yw1NyMfaYbd
JI+YC9QOyIgZ2qv3GxTPmoknNKnasU48sc+cenf7bqVA8q6ATiKN4yzAindFTssZ1qMbBQaSLEGN
w7mUnc/IF2/YQm8CUMF7KNZ6KqhFNm3b5CJ9pGFXb9WLPYsEXsm/TZMLp20iQ92+nYt1F99A107+
/y+5wRkQAneuKL2Q9iYLOCAGmBqB+4lc4MZ6+0Zziq+SbDsal3eVf7+YR4p65q10TA/vaTcuKe6F
8nLHQ8og7MbIPljBM5U4XXZLqI1DrOdEVeggiEmrJZJARjWzs7iF1z1HgMQ5oyO4s33v6ucQivFd
tO1/4OzYF1kVP6jp3+60PX9JJKuzIW02Fg6Xxyal1Vu8W/k4DazNWaDtGkDye9/WUg0XENyj7a1r
6lgXA4cXjkfZgkRbvsJFM6mtJ2O6bjgJU0zmcd4pxi1rH+o+MR2RKdxPJR4yW71nMlDSdXbSPomu
GhLaa+eiPi/P7+ti6lA6s+A4qmESkRvpwG9zNVzg/q0xTxIZkstBUzTEXdAUFn/UVhwPUoHhNJIn
LFugEqxwjfOWbcUlqZmaFK5XWhVG28XFYQhy0oWeFT3/KFR3ApDolGK2Zb4vvpCX0JbbK+2iAzHl
W/wXNpMCmgpHOgdUhHMWBDQWd601hZ/8vKw3Pt69W5Z71ew267to15QXbcm/fh+zYVhLGcvAOVTz
0LLlUFxS991QO3VjW3MuU3Ky/AmM/4zRO0FiERKBLAyILlN7yRPcGEaXb+eUuF3iMXrRTEVJLT1l
zGGgmSUH48YTFdt1HRGpmOUwKS11THte4UHbnyUAvPvmcnkKgGVcjHQkekvlFdusmySF6YrqCuO6
tRYUzWfksGJH0R9uQM5yB+MTYLWzh48FvRrdKKwmk8+0+g2wrD37OBj9/uPeKtdOIc/z+ldAdlwY
eexAglfZGD4p+G4QQYwu81iJ96PRFZtDANcWt7r52JXj2YnfKVTv1O4YGEPmi6MvNkhigY/8MpML
pJkQd6PqLgCKU1OVQpKLgrc3z8hmHrBOCc4YC2pg1jiFxcL0d8CaQbY+8pLQDjzI9leGwyG5hiRK
DInSHtF5wbyd8SRxbPuPh/n8Vg+wqXmJ21Mve3dMubEtm+I5u2bLbZqSrwDMso1/cZSV51NvHZq/
CgCb4FN0HUyOFwYiPUao4KTLjY5wniOC+FOLMQaOGQSh3HXq5zbR9PeAbhMHnNAD4ytdkg70BffD
ZycajQ+C1w/i4sF5htbNPNpgT6yoJAVGq+k5VTa0r6lrLIsVEZ6Zp98z5+8EsXdrxzsd1Ll2L4sN
v1BE8shnaJmiINn948RlUY17aVe166uH13TUN3tuq6/b2csKSJvvKjMWJjtkmvooMEIk+awYtqc5
rRCFXPa2p1SwnucEcnso8nwZscKAbZSTZ/LSTMn5KWs2DzRwSUY2H9kVxfXskkPdb/s3JMPbEGtI
fk00D48eLX/PIhd+caezw411bH/xEo0fXQcYMjYAOILwlwKEyaPvuIqJorns6niFpyr6n4UZEy9P
W7DaTQVw0aYay/KYg4CVW6T167KOZtwMQRLmvJlKu6aWJXOoNazEIS2x47o6Mic5XTBXvvfgHhm/
x3FARe9t8umLwzzZm3yFNYrNw73S44fHCuaeWp6hc9kqLK/s+R480vurRi+eVMnAkpLo/3ACAmRS
3rDbZI3sbYlm++9b3nT3uFOxzYnaxXlZEKu8OS8Zmq0ou7LSgWT0F6KIv59VmEV2tS4DXCvp5l5i
ls7rPIxMkQsn1ENp/CYMEjajipPNKpjvH/UfAhqicMrOJcUBkU9pOlIBDsoLPKEqqEED14SFYi4j
YwdHshtR/KyA42bM/g8ebTwdRi6aj5ASmQzSDX0DhN+muDU97emwdXiEQgVBl0Rv5JetoHNeEm+E
Bmscjl5V7FAtBJfdzZntjOjhxIRWi6gqsJhBLVRWIfr4YaAIDAAz3L5CIa0qh6ci6F5vn1bEi/Ni
3GDMItpP0a7FtSiBRTnOrtQF4nEEV2pgHId/h0aJAmvi4CvTrADp+nqY2zbug14wFaNgX6wI+ltA
mtBW1W/s8ZNuROgKejkV2oJiApoHUpm0oDRH7M2C/W3yeHAJzZpzxy64HDQ2GMPuwkBLBWJS/3dX
1OziabiIGDfP+9TZwHzKCvyOHFFPW6TyGhnV/wfDdO7SM8c/RXApgtRMGVgt1cK3Ke/PyFrLKanV
SPhUlKpsdsUsz/Zuz82WHbAkXYuKtlTjMn3itYBlmoYu1IUEysnpEPv5dzLK7ySBVKyMrOHo0DUX
eIjzPJuhHXOEo5E4hXFwWx+2RXqlmKomgdzcpL3PzBVrTlGqn6uUhrg2JnlkCKGVTdvBCiN7KVmD
gRVudpGj2niklUIkhmJU2DpKrjhc8TbegXQWwQVMMR69myoVrZ+J1L03p54NyfsimGj4iKebnGzP
YXeo+27x528jgbKWDToNeHHt8pkicbk0tORhKz7IJ4Mxb7YImchvsKF+kp2jC+Z/pgczpkNgNJMx
lRzwjQb4yz6gs0gl7dmaiQBkOobCy44e0svqGWMO76mpXzvVr22Le/rAP2yxi4qM8GevzP4L1sJR
YsGFvUnYruM/Uw81BFv2Qm5a2konAJl4xHhrAnZq+TKK9PixkM5xXdyMj1vrFwhZZ31fwCKFWKHC
nWyC15MPEIBDk7xhtDN599KDQk9U4He4UnTnJnedbDyiMTOAUHbmdr0tRpKbDaDOcIG/I0Xz61PJ
wEKzE+WrmbMU0XTX1yvlIIX56VKPvTEhrpOFciNPSW3XoFHaseRt85LjzlSJRCrEGlrPCr1TyTnU
F/r9hNdgoVoAL57M3iH+qYRNLvpE6pAMWxQadTouceRpxtGoytWobCK8/17dNoFPYH+dDVS7kwtK
IetCHmVgjVxwn4vsnAPiMBET1V0hV4XQGNcY8nCbfhQEv1QKj4+wxMVaT5xPZLmvf1Ni4dSgECoS
UzOPyWInpfq3QkYX4evx5DJUsEm/ct53EMsqYkFeLymkwVhl1Q/+skzbFQQjtrXIAf+y8/AnsorW
7fkVPerNMWcqgFOuZ8nY/46CIQsdaf82iYXayJE+7ydrB4vh6nmujl2vhDma2ee2Wts5al/xsHOm
av05umFXA298RfPDh974GJNDIKKEEGiywa0PsJrGEBGyj+Gr0JjG5DH0bn9DRkG5gQhPg07Uu3Q4
n9kacXYBMBX4tgPSUTuDC5KtX6DfAPkhszUDsYa1+tv4IviTTcOMVLOAavaToeXcmWRnjn2B9UMt
cdscICgB6OGUnswYpWepY8Mphln4qZqMAijIvTKWTn+WVSosiHdJUKPuPk7dhUanrLDgw/fOX54/
Rhawus5jz8TSHO9sF+CtGvOUSdHNakFhK5OP0ykr0peOEehP1NhC7gohH5hzZxjiz2lq9WEZAMwD
BeMtOKrZC4jjxzJr9/xzrUTm0/KVV7WZPZld0BUxA9pfbueXMXqLT8/XRLSUCGxbuAChdYASdZ5W
CFvpv7jFpQR4jNbPDtBDxSpAW4IzZgZCVMbe89QH32ANUeHa3bBkDrpsUQi5IaIz8xmRZuhtUf8S
PlzgBhDfgS73WNT1RCTkp44tt1EZ2X2HNRKgIZbL17YXxfdQRZ+0hkZJMD+Hr/63Xvn611trkcZd
PptwaS7MXzwfiIIadfMKZvBDGcONR3warDHbzTw7PxnWPGHdAR6hHiVcEcxlTo39OE+EPNPL1vkY
yVJMErvLnOwFDUWAe0NBbSSIMOdFWKImRSX3DjKH9pw/cFriS97Fi3ZCeN74C3Mx4YCCBIcHOf4i
nz3k6B1nBv+1ncpILbUASr8108yOLJWSk5+W5l5+MbvloTyfH7jdG5wPwpCB/Jfod0YfAOUYiF71
StsDwudh9Uqkjh43RklyPpGJemJfM2QF80W25ptbLiTg5aXsU+V7d+aP3wqRIbTgK0N9sMDXNctP
wiY0VjZxqencnzSUW8HbD/+/NrKBJrhUMv11Y5BAu+hTknAgUMDm4/V9C524JfEJYrpa6swGrRW6
5a7SG/dN/mVZ0mrwLHntHsQb+gXZMP5rkk//AeQ1YRaTQS8z94W79ImMlKJc3a3GFZV/t5MhIyin
yGa1J/2c6SFtABKSplKXOrB7jQu2z6aBa3RSGwlzHg+j1Qa9mbqTGV0t5kuR6/0AjO3k6TaShZ41
F4dNcgmdA/9UUmPUtAVlD1FWkH/aNLRTK/XVexnF7fplA87qqwtX3pmT158E9QBjOhHY+i8Qcyb7
bm205ImCoVkt0qoKnTgdkJmrlgaL/E7xvdJxv5IRdJuCsFBtl8/7NdiqXMwwS3SV9yr3sRGQVvqK
Yi5Ae5cP7FSvmdY8baGSH/AYicCUERUNRfpUseZmRsjd2vRvcg4Lsst8Smv9wEe7uejN/Vj9Bveo
xTX840t9WqJy5bPI3uPP2SMPqIWgz/ydNvCPF+cmGe1sagX1f4rApFmuq+0ka1SX/Zr4jrJ/nMUs
CV0THLyoM2M/YXtVpYLVhX3WHUXKVL/7rgrqoVb7Vk825AaN9MkJGHpof8WuEsA8Q/bEa4CrikWE
lU+1lC8NMaJh0JFX40qeLUhgGkv3ZkAV9Ql0Ydf+sfu4V1FMw+DgF5NeNl5r8XhXcKDCufaPCXBR
oPKnYBWqghoPUYXD3ELnpYjJnPVNiFdNsJx+sNl6Z9nOYxyYNgliKvXK3YNVt2Zk7i4HVYUfJxPx
pCYUcUx9N+tNJS7TolrVCvVR52vx0vQ3qgyt0sPg43EjNeQxV8S9aBVK5bUM1u3f3Wuur36IlV0X
DGStEW59IEBtcrDQOP/TLPrZTWBIbirBSi/5clHZYrQvcrkS9MNCvnT0BHFUWBwFzLkusZfhDVzL
YdWwF+LUcJM6M78XqY8XKBOLmz1erp0VjN8JBzDRw6YIJgAgI6CtjeVIuvP/S5tPMLWwxGHXKcjZ
GJxYulcVpZTD2NhD2WmATHVpPnIMRupb9koIXxdf9sCa5KPapM5Q72avgbSG/lxDMleay6aCDDip
aOJJB72DmPSQZyC/CnQ2C2bVxjAj7TnAtAk157MzqC9um14TP3itFmO83modsv0AoMRu5KBIrz2Z
SzCPXYwDEGUQ+Rbz5MUK9ThmtqGHpBdBO44csaIFRuGdH5SzCKlVNHWZ5XaZVp2yD69VB3jswYaM
hck2qnDMES3ieXVxlv/alDioWoLmTaDTqmx+Y25GPSGKTUSshyJaTHqW5pCxNG9J1OrC1EgmvM4t
/2Xgvx58T819ZVQ5kBwLUgyiRMMgfIZB2RofXDlX4H8VdJdDqBDQpjirn19cIPYLQ4HUJwYBH6n+
nnJRAHQB9As0sS5EOIe0JQExf9Lt4YdvGFOGhPSYwcfRZ2xDaatpnUhfK/oAUKg5NT1CZKQejYQG
y5x6byDQan2fuP3SOa8XLH773Gyhv8uQSOegioRaCxLsjqzdPvCPBoCohYLwahZZz0L1S14OfVze
vwXuCmnw6X9zkuCB+0qxX3PSm1IX49CpHyazUZcRlo12g8fvFgAGGn42Ae28dhSkOF06LxjE+YfQ
kgdPPVYed3+XcYdL0l6YEH5V2dPUqiKa7OUXPNPyj0/Vv8/VcKHiUpT8kezkDj4KJAv5inh++13E
jDmz2nktrT1FpVq2WraXHTKVj0yGjrI88IokWOjd4th9ODG9+ChNJASvuJ9CEWARkbXSamNd7TZH
a1/nW4X2ccL0sOrKrYmYw5POdz6ljD6um89otG/vd7LriAC+0iVZHe4/A/4EpefR3ZG3LKH+wG9e
R7kUbsMkOwj2wpQOCbl6j2tf8XEnB7po1uEmyYQWuu8FR6pPqBOKzF9YbXVgl4omIlNJ3uQc6UW5
K/RnxOOv3oIXI6uJrFS4hEq2peFGUTabcd5UgcIe9UD9O++IwAqKw16QdwbByM9BR8NvTCY7GE5p
c6D+PBapTXLlyskwqEFc4QLKwssXkZfcfvGSHBc+rV6/x1PoUd1L3AjdrLaNiWSGG92Kou174UN7
o27BTF3kbaN4tOS8PFmbQtysebtzQONNl2qSxIL5AJQOY+jhl5XkkK9rVI0UuIcxvxU34m8TZRLD
ETGEF+zUGPxX0+5qMq+4XcZ/9/WWWOAkXtQX/Ue+8iTEX9gD4uJDXKULxjiyUPgXhchSHvfz2LxW
DJ0m6al5CqKHHhbLy2xZuTSCgvhiOQ1b3eytPDZv/R6jJD/2nbmAQssbMu+D1Ld4CisU80K5ntUF
pBTMYUjG+dE+TilISPLUK8C+Oc+oaGDmEQg5pPjLYlBJOh4LWPPCH8BsdExAvja3jDm9y9ACgo0c
iki0Bb2rpUNUkY/KWqoac2+yBSjFndxPDmy2hLwRmTHM0EkVl7oAf9Hyaw9J4SQubqbyLb1XaGIe
uDwJTPC3ckG/SYx2ntjezzTPHRCJqkHPnsfh2HFXoBUw2MP6isfgEUh2aU51yyqdnsOulz3eqjrm
sUG5hUYeXOVrAzqv3nxXLZgDwanq3zYJJRWjK1LHDKeEHRdTcY4K+Q4E8uMDYaDtoTJJPKWTbI7f
IwsXPvQWBp9gUrSyKY0LeUMg7P97yhLzvIIzodvz9jpN94lACKUxfePfK3NOLkj65Pedae2lMsju
g7jFbsOwgeY2iIwUgWH81X50oKliMJKhNcS5zyu6Zyz9gYHHnuMagnGjTUb37XHfenTiRM6tYecb
9Ci0N8S4zqgEeT1J5CcbSVOpGNtzDlcjawM8lTBkijZqMAJxTqHBqx/7DIOAgV8/AY44nH4y/KOj
NWQHZbpjzc8j+VlWjcC7N68ZvWPCaXXIFXWmekODfGTK4lgLCpodOprCuADRgAZlHOzdLrturNLr
ucVMDbXIlK/Y2lnUadcgYaoT4+5+JjU80NYTi3EV3pm4lpNJaNUQtF5gYkH6k9Pq6ex4LjPgEbFt
IeJdk0axLQBwcHGeaIIF513Xl/Z996xwg6TsQeza0DkQaVhnSKWmdSxnCtdoFwXRpgcO9uH721Nu
X9EmgEGhw2TQ1134xBNrJ1uo2BrtYH+KyfhLQLZ0+4nSRbQlQEl172a8mPuzg3MePOYIKQlXIr9Y
nC3AOVT9TNOtvDG/JUftAnlpaMZ7sp1pIt9kqRW1iQQOm18xXwfwA7zEbA2BULY5/xErQYrBl7fI
/4lcw82PqXzBcitQud22uQwOXPJ2Ebr1+HuHDxnX7mkFhwa9YsjKgKfW9tIcCqOENKqVLN0Ch82C
PdqkfqEzz0lyxJM9wdyHxq1sMLkQk3FQQV7M66OviqQxmEoy4NSa/s+5qGX+MaQ8zpluzGRFlsYR
FNNqQJ/Xecmqc5OvChmMHNTWF3spTaGsWVhpHhMLManYAXWmI47m32+AonRUx6OKxl7ahQW7aQ59
mjzqv57mqD5BN1OrmSth69z9Xc2xAHvDbCL2KXaGj7NQCd19QSLn0kXlKfqwVYjdFrDR28BNWCdv
UWKN7Gb5lf3RqCAqLRkkYfVsJD+tkZG9X2eM2dh0joQ2jk7880zob6ngxODJKkYp7ZhliM1gmvq6
KZTPpp+53DaUj207unzyFfZXF00+wMIv2U8EYmxjvB66siul+RtYGJqUeLal7XJybCtLRU6YfT9H
zNCzPLoRu9OFVeErUkEV2V+lt48KpoFYOwh6JzRwGgf8Tos7CGY6zL5I1BrGbRz2S1mlXh4dGKr+
liw/6hOIhST/M1f+scBDTkINMy4wKBJfyGsDSTGOhfMWxErWQbYI6hZFhrc9f5scl9KGV5zrOlNV
Xd26v9xbIaMcFCJkQk8Rs1Pnfj/PIoWNoJDNp2qQxMsJvXOIMdIJpblcaI64362TzLtL3OR6jQza
Jt8hdcalvbl+RW7laZQwFNkqMn8JWRjNGgbKfRnF+14eg+Wjp4Nvqkz+RLz+A390YDuFxwWPR8t4
JwdpQB+vES3s7W0LPkX+J9dVoRf9zpEXTjFFaA31OXvMXLJqCHkFWgUGXcUMO7bS3pEi1rx+NGCv
1DYeXtwdtvaZXoPrxj1R2ApS5ScjCGDrqXdO7r3q2vtLrtfqkjolnYE22PrlmY5QYxqJYkCTPOzr
Qk8OqUAQcW/PXy1AJAYttZ/+KItbu3tBWunZnmw8XRqlPwBr/uTt7qK/EpP63RBKzNFrH29bsUDl
iH1TiG52t8XUblI1mw7UOEQzW0DOzQ7jRDW9VOGNwAyGIXuYhIoVx/p/+gGEG5ZRfPfO3a55dIXX
LWWUGsWqegpreUJV6QOesIKqqJPGTJqzM2TccWHHZt+2Xe6ldXAVSE2Tl/id8CNjzowhnm09Je98
GUlsLKuFJQLNOTIlgr9t7xA2sGSYNhFzq3ikcH+kZQaYPDTIPXR8chh8iZYlJA1Wxu80bLTFaa8i
G6GuRbvRsKxhC2Erp67ch28x56x0dSG/4WaBnudFOzsSciFMqEDy46s56SWmkH5yiJKlYjfU7IqH
3twZoZKrN7em8hfHtLmnJAm2MaESjy0OmkEUwxbcAxZnCm2lvHmpubT4MqJXW9gkdibm54iQrUF5
WxtaAB5TpeUqb25kIAvVa9J45qj7VBDMn5jdZiYKRGmSL7A16NLgDC0MsGG8i/cj4QcjU8ptxz6Q
FzuylEiCmwPvsjmVG08yQ2tlO0U6yiineFxF43clP/tvDXUEOGeTYP6ZQeVq+TmAS2p6iLDEY5+s
QFwZbdiJzkLWizItG1QoU1jyu1h6oRyqzDYNC3/p95CDx0N1D7Wo8EuIgdYCxdzRH3wh5FwZg+H1
1wUc9H15ZqGiPAktRJv/kXGcgY2e/hlZU2FqfgaE4b6zUjeZnLcXiRkcoVDbMtHIFZ9Po0ms3XZp
BF0U7vQRS4lcgHuTxlvhJ+PeJD4DB2VgMpvMdXQvXqpluqEeEK02jc0RG8KeF0o1KlXwiZA6f8te
ZQoEpIGXTVWKU+Q3ViDDgXbjMIGxwpjVbqXz7fc5l8hQh1h8UR5K7epT32iP7/c3nCgZoH4VIeS6
GyMltu7SaXzYd5MiyUNGNdVpzjkbwZfQDNrPj23taOYRzJReAUoJwRjWutpegcDFO1h5Cv2p6qwa
qbTg/vnK0JhjN9+Ogr/BZNk7qyLe5JdLeqmvqzmWL7x/+jtnMdXZWsd6tPHKwJlUL9fXRiqluVZF
aCznfzD2vSD2mN8wXGVGPdMQCX0P9UdiXXjfQCmJOgUL+6Yjo6ABLqFPauswR83N2N/MaYDkoxZj
OX5Nax5Ahqz6OIUdBWYb7Trd/whajRDzLIEXrmT90WggGMoRCC8mctVPHH8sL79mzrLAkbG7Gsyf
jsjiBbrSHYGHb1JrQaQ7R31qkj+eDMN40blFjmSTMPvpyEJ0URmJ6Bw13+xmA+/7mmZk3AGKZbro
X47DSF4bDh6G9MzzLE6YUO3uAINOHejGPtJQxOS/KAIkQ/+Avk1iPwQPwiL5lOe4+o39ilFnLtCV
EnQ1PSKLM59y08CKrGwrvnRoEwoO0ONee3bLomlaVV9VU87NyO7I54caYTztkuUcYfVaubKI3l5T
r80dEXBlKoX6CLukUZnQB/+R/qQF/5j0n5yrCCVQfd775ZMYqMDbohxrmoQYCTisw/QS17dTdGAw
5r7pIBFcKEN7F1pzZqHfC9Kf/L3hCRQTP7H1oi//lsKqBNcXO2Ity41aXf27qdrJtJSuA70EBBuM
d+wjGdsclpEyVBOjtZyd8uEglyHh6OdhQUzlhgCLNsFnq52AlWEY3QjHb/+UgapE0WPwLzPDxtIa
0HE8QA319h7bQlAaVwQpiDyCR1DdHyaIkrh6KHrcL9QK/NFYm4np6Wdx7VkJLVEBePNBf7YmuR1n
7kPlrjYJIYirkDhEP2tbVyJ6BhzzgVz5bnAjjxsnBqAbIrqyz0EmcMvyfOySkUQY4+BOiLiUEtQh
9zLc4HZPUA8AwQ8suBcvicaPWwiciUgHDdtxoCkyvINUHYzoUusN2uTmxTwqYulswEPrhrJbYvTt
PQW98RPiF+fI4HI7NkWWY2Qttic1PUPKmgj6O8vsQFLqXRjpqOFYhSGNxaI/pH2XKemqrL1V+BbT
vZ+D5WVGBu06aeQQ2/3GCTtxpS3+QWHs2I4TU1c2lH1RFXgipuxrQ4HCj8URJWh/72L6RRDREzE7
AX6E8ByQARAImCVOfrSpNIOkucdEgF4pGS8BY4Y3gGRPqd5oengo2nFSpiNQnAXB7JMi9tMK1Hn/
BydC5WANF7yF9y9hpdFaZBNb9IvERGZ0ofVl2UQ9q9ntJ4f25ugbqzThlf5v3xFw1dY15vEh+ptB
DYk4DupwnNcvMwqqzjSBe54AajT67wIaJQiITAtzCRxBTkspscKDfiUD9IOWpTTAxccwAv/oxZFg
Op87zQBh+mZtqqhBxG0cM/uXzmC4BjqR+4xVWO8knxxlG2SgFZ7FZ16mbbFzAkkyJgH6PQv3nJsE
7VJUTtVMyBBxJxquOQU0+LH3GX66CCv3aDo7sAlQcP+GC/n6co1HxJE6ArLdP4L6wr8VFUX6zHpV
9Mf02KaU38zP0qCMDd0gDOexy4OcXfTaQPzNbjTKhgAiBSRF6Yo9SnQX+5w5jSxs8ZByPNtsjlpj
HraMUR/uE6gMh+EfD1RJcJr0oQJf0qbkdR6EbSX9QPy0KqPHCZJkKF/A0hYQtOLb4bSmLWMt4k0y
fHiAiV2DqwzlwG1gAOPk5HWjgV+PkzhJHFZ/TB3y9UyL6tXa+OXZApwE94zi5TtGSpKtihCRUex7
qHRTwYEQjLAxwlR5IXwKgwPHtfInjSgD0pHZbDORD8bTpbb0fTZ82TJ6CZX62jE621acq6t4FAc6
p2nyTuNTRLgRz1pSGrKfRFC3a56cnM+tBteG5RzfX/Sh+SN17SdWDdOXSquWlgDVwebmpm05cefi
UHffeEI+19HObgZsgbfCWwQHJantlG9M/550aFlCJp7Ntwwh5avDycbhCqkvkJqEVKY/23N2J4pr
wE48Evc87kWOwM4eEhkyZYf4+IydQYCWlluu0WPcd7maioEyWW3IpoEs4yFoUHAoY5oBAyy4D1es
A8VU0HvmNnMMWZnYuBbPb8jGVnSgQhIPEFHjlI3Pjios5xElXWpC6abdmaQZ8uzgvUUG+4fFSSpQ
9OeTuluNts1wP5rAFTF9K0bxUbz+HahdG5vsn9eo/Y2/kci8kLhCskqhpZL4LNJ7fC66zPTCi65E
dsmFa4fyRUxOD/WGiRy8L7AdBIUPVAnLDpCHZKlHKWc7y1wxktJMZ+lGTIihDgPZAqy8YHzqCyke
7P5/5G0ODm7R78sTEOugCKp+Tde+lCehKqQ6nJDz9+NtWlp7JnyhwO4TB4R5CgDh5N8z/EJfAnpS
kAxikBdpDbJOT4NvaLryEkh1jr1Vc5pid2/jXFvispGUqsZ7bm9kdUgrO284WsjSBsxIx5VIs8zK
rZ3QUOc3TUVeUZj/kIZ5FBRM8Kews0J/SwQkGizXyzt9rmrwcrYCK14FFZiHW2P8jjrv/sx7e8P2
2mntOVmgAWCJoI5exEsSgBgrBjfvE4SFHfUuLVjs47A+HmgRo30FlifLiQyfz79SLihPEFsBIcDE
GB+ihGwD8GJLhgcZfkFaf4DiavT1DDWctVfdT6+e92EGDRldGMZ7TIRyW+K8IVJdNTAHLpM3HJOn
/g1uK1Qjko+umwt0qubU/qY1BeaNrnZNfmSAjwvnJHbyIqcx7Xuq+IqIXsD1iFYZF/SBSeomTuIz
tmGasGHSnpQjFsfA/EHsL2p0q5QnBtr63DNMP4ao+bxTdDmYXQL2mR0YIzn/jXsZNanmggMd5oF7
USvTdtabePQRYfoQ/0plVOlP7CxFlqdfP95TJwrF+naXjQLAeiJVmfDSgOoT53m3f1Jc3j2eWjhp
HCBg9PRRVlg50LcGC4zJiWPJgoj9jO+cOTQ4KLFOu8QVIHl3OluoOp52UWuoMXNe70Getej2+g2y
RQ4AwMr1WyzJIKrZ6P2U3RyxieTiH/Nht9yHtuNie9L3cP5QIJyRNikKNcQq5U7XkUoQjHZ8t5aM
+fuAmxvKxIPl3u7ZYUlfOFqskxYX45lYsFSE9k1JBvuiyOtF7l/TNM7MfaGXPT3pCnQ1yHwzZCFL
lIig46gXVK7mqONHj0D/veHAiG6cUcQ92WsHHanPWWeLTLAv7qaiFnFuizV+KLRUxOTe9U6vIzkM
llp1ncsk2dvuVjIhoQhQvsT60e6BYpEwclDhUWG8KjtO54zUUyQWQsRbF+1i+D+V1m+FrHTRyD6P
X1BP6YIekTlhudG5EP4nApXFB0Sx8T6VGWgKN4JXROX5hlZCzl11nH/j4C/afoelvyDKiqDfTyqr
tn/EcSQwX13bXxKDvM0eaXD4++5Dp9pzSDvD4sYF3QyjauT2AdyQdBdc7y0iUUxQ6ScBZ6wklQ6T
Tgeo0lK+flIO5OrBifGcT3a0wdpfAOZQeTl65Eh2O0KZJ8c9NReq25lb1plyeUio47Z+8kKaLsWo
ikLnPElbeXc3imzvX5dnqq8kmSD6zzgyU8+gEwLmERRq7OLCm2CYSBiQRIcMXj/NqhVRJ3nKYs2/
eGVjmheTpfldtp4/4wDOrB9HVqidBRcu4Q/r+uZxYm5ZEO90mHFvccDbTEgOztZ8KMoreb7cR6IE
1h/cCbwonu35nMZutSz+CQma3Z/a3oo46Fj3ufBlg/DrPDWQ57g2yyni/5q1lQzpEJDIstlf7pya
q7Rws0rrrYYFxQlNWBRUGA2oxGPbQ9XpTisN3Gen78W4Jnsj2/qrVshic3/w91CIcQ3SOyExnXzC
AKxGcnoItQoGT4h0BDWxs+1u0tU0m8CXGTmPLOcj8f8H/yyZoU+7oJudJHnCJ8AggmC+U3tjQCC3
l9YT4vIJIds7U0L/eI+BGo74Jcz3T2oxMAsTlfuYLZFcFuVh+ZkcxIgabbGBWVz4XdbSv6zx6AOT
12G/343b3CHcoKz1ihYcbwGtZVOtgPw9skh25VcfJbMeIuHZxh5Ir+ns0xMcFuU4qU0eC8Z01jbQ
vWa/KzzZZiy96VRefHDPOJgoP/wZEQINmB7TVHe9Q04LktT1SWmaRPcV7U3m/LmSUXGDcujUeb/+
PfQl4gmmXe3xUIsUFt5Vo66Rh30qBItfVKFLeo1W6gZfsZcQBz8ttiBHi8gu/CGPNCP3GEn5aZpY
RpLTxk0e1YGAhqNF7evcg6MaL4ScmgJDo9kgNul+9njYH5/y6SoxRK8RM7MEcYOKFG0AilurICKv
3kP21QidHxVzcUpLvdwACk3tXliXA9mcMbFaDyx2rVPB89R/nU2lZ2cN5BOla+LWF+VSTNE5NAAQ
NoVFeei930FoEbeK5N9gxu70Zu8doKtCXDQkGNv/DXh9ALC9GShgyuME0xHDBAyQHz1JosIAA0u1
spVHrBPEkXf5/5mH5MudF2jK4ddxG1EVlxSKS5i5nRgbshaQG2n7z/jzCPWU7HJyILNQ3s+sk8ag
pl7ueg4p1MtJSt9Jer8Mw5Mrdochd9qjCVDjiRoHmjcihUrIKDldKaNYgxvCwQjDajX9I5f5N/jT
ImOy6PzXL+g1ml+oPgLh/0syenOnAVyyDra1LWJDiV6t1rsN4NzJSzGQEFk2N9kX78Ot7eeM8ihB
tU/nj0FzDDj+2crdW5aVsZ0Z67KrhQFZ/S1zQDfTO2pWLLANeR1Bp6BKk/DpAlqBLoTXer3aBuZe
bmgXaMjaTnUC/sXq0NNcSJmmT01H/c78etGD0lHicQHnZOxRrpDXA7c36XCdpCUO2K74eutRvE5v
QNtjg+JNC3lrauOCEO6WzfMvv8aKaxYBihLOPIybH4lONL46EC8ePWx4+VT1sx8Q6BzhZVy05YXw
hzxTkAMuEKVHVajuTnWqPj0G99Il5Iyzx7WsM7dAQ2fNoA0FvOtGF7g4U2zXb5cBT8lGrTBN9Gyz
ivETa2kKOtiIYnUbFcq2ashCvGw7NOVIV/2/ngaM/On8rBaQUEMK4HJUgrGQ6jPDF4WM4Ir8eF0R
PBItdFSYO0r2lK9pCl+YkLHhGk5zvnkvcahmIcj2TBJ4EcG9fYgsciXeYq/RAIbs4TrgjV2Htl6z
+9RNtAkShoF+AZ0nV4Bz5Ab6RCw1qvof+lQ87mRyLJpMZjq1NiuO2In1mqY0tF3gOMzqrB1Yi2Zd
IZI4u+O3AXfvuspSMB9GXpe4t6brnrNNJw1QVhaZSoGEWH0Bh8ABfkPSpAZBtt2G6jQe/7FNKCYV
mIJmvl3VTM547KMtCwIcfzJLQ2OhRwQ4n7S+FOJXmHWfX9n+46U8QHNOctH/1NsUIJEkir2tI96l
+4VRt/w4QVssQTgYKLi9jsai3MgsK2pcFeqxyomxsVxdt7VZXkeUEIWFFRZop3bAoetDeYw76K98
riHMsm+UqKCGkZ7MlOdygETb3eDbovSu28HTTGmrnmclQTrdCzMwt5AoOFTy67IPjMUVS5x2Zi+D
b1TkhzAUStzLYHEYO/yBHRAG6TkzQ51ic80fhG4GikZIt54+2ym5rCKuDjH8Lh8ozShO0419Zq7I
l4AgEjCS4xiJZ/aljg/qHSXY9L7eKVJXMaRK9meAXwXd0Fd9aIHQlsuWm1iJuS3BQWFIboEHtQvU
S0E5NUetQRWfHeLtDLQiZdb0D1rrrfq/XihvVJWicrAq6vtSOZNw/E8wfQ/KE7kPlh1wwa05EZYv
gUhrLbxEbv9yKam430AvmzWVcs1qUi0UQHWBQm5eMJnobAvJUgNy1XV7NtrYHPGgGApB2px/rfNA
xup2bBhngxWCBPenQIAACe73Nn67CDHm9yTIHVZY99OTSOoy/vYRC1eUISMF52Vgv8URQprjEE5E
XoDPCJ4CekSeS3XW4y4WKyDu60yLdFm2AcJMqQT7lSM1btOYcpV5C8EhwlFjLSXgl03/jhkfLAkK
Uyala1tFv91wtYmMZIZnzHYqb8x7XSXSnk2Hbhm517kgwMSV1lk8EOYD+XntH+VFfh0iyQ2J8Pip
f+HuU4GGvx0nDkbzZYb04rm721G9CtXWjnxeRPTbyRx+26Gbo0ngthteBLOKQyDKuziwGhDVL9EC
yhBrY55XzMIjo+NTC4Tb2HCn/eRPCvTyspn1nbKm0+tsC3kTkoQmnw/ZrWFIugc/2AkiQYixm0DM
y+dm4uiMd48/1EjuD73xlJWQQnoGKItEZP+sAVAoVnrZXyM9kWZJRO3sg0YXB8Ca8YVSazvDfoTo
KPbF4Hv6Y8UeRQ/atsRUH2U1PkFq1lZtHuxWi/SY8ig9eq5ywoR8SAJ/yhZ8QXxIy9+RDs9327As
8fsKN4wdUePMB2uAmedoVR/WY2nM00ijGU5pRBdd/3IuGWG0LMGBAHy0Iz620vRahJGz6DSwZSkt
wEXkVvxXXAuIhdNfbu3D+IpSFLJrDUMbvKWMC0YbJsvl1ErdGbhgY+7Bc27QGlBEadPGefpYAUV3
ICkXZqAdpSmuI+Xyd5K2Q7LWDaMlEW+gh16VazRLbXiFwW/oNufSj9+g/v7/vlJ2kNmr1Knca0zw
XLDQs3GwZueju4qok2P4DnaUHh5x6/nfXhItQRGXGJetZzpQ5SXI3p4g6GMQBLqKoZ2onv6TpWx7
r8t25dENWBeIbgUdBI1WO0S252KmMRa3kN9qAhoYezz6c7lyQieAMOEEuYFaQ3zYukzABCnpGh90
ttf0w1OqNlLGv1xxyUE9y9Pz5YfMBEBCLksZ/yuxzyl+u+ikYLBtOfnz1hq20Iz/NYORKd/hNJST
kTU7uHBmZ2tQ/qO0giZIhwrXIDugPCwFS+UYR+LwWzN351DZZE0LnveUoYyupJy+MT7xLJbaZR3G
U4h3hCYGVVMCX7ukGCDcfF6l8KQmy1QC4AdMAXgpqm25O2/p1RTLstzVqYAm2kv+KnjZl7fA/lXW
44gp1sgo9njgYUn/MGd++4n4Nc5E9tNianZgl5HhHI6cuWPnHMihLi737GU9tTkI19MEAfCfF/Ff
ePc98oJMTP10+7V9z+u58fvdZCioofxaq6XwWWUYenuR9dRGg9RUfi52oq2S1Jwd/oIxD9Xd1S4t
Sau6ITPus5YVO006EwEU2iyEHaUxlPycqmiSwQX9Ayk44hrq5KeHBSnCd7KqBYyP5LgVpf254GJZ
Kadm20f78WSawoBcOTtOtBCVWItg9v+d77TDbMOI1scooKqThPvoveumei3z7g8i6X2+I3GL5cNk
jxYYLzIyf7D2abthVczSaVwI4H819ujyShGnajey0w21ictoq7JhrOv1gwiPsRx1to3jVk6H5gT8
b5z29FvIL+Hwib5cs3X3PNfOyNUVsoukm9PRMXJSeUgH9lEvBL8YF3hS4myvAcJESHR+uCgDhKXb
CTHlglRh6mcOGYwywtoZrIinmHUaEFSXYEKEHXZuvFJgvI1GCBa26IxWJaOfURjCvEdGD2Tnp4ao
hT4kw7AzcOjCR2vWmdx8yw8fW8uYjMIryx4jWqUawuaT3n/cNJtGX1NY0448sGf1aL0R9Hf73gXf
XRIgun8cMkzXTSUdXQKXUj6qv94s8aUZ44JEeHkfX3lSYkmW5UbJqW0P2srq1iaJ9iX2eZrdF6zx
GcZBWCDip4y6wRY8XSnplGG29gA5hxFKLRLrpYri2JAzaH2C67Noqw9IuvgKnQuDf1/jPtRMZU9a
USZPgH4AMxD1ilMKRqpgSq0UXKJMN+8eXqxmqIcVhARlP847AAShcECldJNxxpv2y9HGtwvhiO8Y
eATC6v7j0N3+v6ar+LGRRI81gRksPQS/SbkHwdAxxzOuvZ2QXnjAa2vFkC3441GQ5hMj13af4RmO
HCUp075DgCO24fXXR81dHqDROlLLsJp7BNpnCx5pZq5KLETUchKifzJ3XY16gKrigtxhomR5tTRd
iG6cDpZhKac8RGx9cxhfI7qAxZjUreIxNd4SGYAzx8EPuHNiP/2LQweqqOFVBflOPgDE4Kt+5V4C
VxO1fDz1rGlaQ83YrykNF7Jxm01jSetvN+YT94UbTeJ/4kC77bPe/j8CfwBFIydsfau8vhjzHWNJ
GbGumhA8xz6NgkurGud8cBODAu9uLxLO2smY7nqVIMOJXXw1p5LV8DnxnLy/1UQuwH2RArFLpQxI
Wq/VLwTxUWtAilYqvxef9yzwp7RkZCCz8uzOwDdJ4xHch7s53McYc5G8g6BXfBWE0ryi32TUJTUB
y9McqJGmlZXOSQMmQ3snnb1Of3Xp+iehle+fsFTTpLVgF0xfBrz/7nU5WGE6cflcGSzaEYljnJGq
YZOXVw91TaeIUP9lz+3gcyee0NSskXKdMEI+1Qx+He1QLqNJiyipzm1OQCOY7kC/Ss8qlFJrrr/G
L/m1giYu83z2CckLlU75B35lXasEWG72IluPMrPNZWn+R8bGgI3sR0Cczrx2bgNm3ItY6FVJFbMA
T1lQ+pOwQVJclUCij4EfyEWl1LAi49QbDkormZl9bJr8qzmHshsjQnJsMnkNZJt8x+Eo3PwaMPah
knTtk2kK57JpAWLXZYakLGXrQNg9rf+hJjoaKXUTsc93FsmKjC6V5r2jVBezyxgFrzmqPQLi9TmW
YJq1wJJHSsthKMTgJs+8IJtXSO4pa7pDGOrI2OFTB/OzwsY4f9if/VemHOXnl9RqgpY2TcVPjfLo
+FSNf7eb/PWDigvxQcGu/9lzVexLNPTOJkofeuMgN5USkJ9OITxvbt2wNo5uM1tjSPjRvwMYv1KH
tQMBWKtqxNSJF1C5j3UyT5xntq2bEiihVQjTrmtHDb7xzi5KY+2gezJ+SghyWGIyRN06z2a/IFG4
w4rs7YJPb/63kIMI40vPGsBV6Z2sR8wa96iIfWdzYDAel6MqqbKCth/12EeJwtD/HKXWkWdW3Out
rfhWLW4GE2u/grL82SpA5jW6Mke4XwDv/LcwQElnhCjMDD8TK0XBdDZe4TmLtIitpR4HSkXGgDom
fbL7Qej+Jq1WuDjCTON+8GpQdQDE7FIS7RLYu0Zpf5XnpSPFHIJ8/ESr/uVlfomaNQXdnzp1nFSC
z5GiHL3FUFSr+fedxKfPSpivgq/qR1l6eN83Dus/gmSdbH1uNPo/o45+cNhkpLL3ORii1pneMJaJ
W3Ujv1wGI0R7e6RNldf54WeOhaU9+jC3fsJ1eJOaxTFoBbpumYUnhOxBspPqxi/pOBarV11Cx+7V
oVZLIkG1ApSH3O7qwuMGbQK9WkxYXw1IIP/zlI0UGT9kOMnGnFENbyMSexBWZfdaXizjQi4VqAdD
CA+TLzHEPS0+Hkr5UI9vb2EIHrm5QVq1BT+2ir6+KNtD/Zx4Imrrk0p3X0vYd23KKK3L8N8qO+mH
FzGabaJbms4uBjhdR/BISXlhcEDgQuQvWVjVZeKggXN0t/xO4Xz+JH8xXFC6Dk8OQ/sNYlp8nUQU
0EYsGFQCEhd9wKsTWB98krnq/J6KRwO6TYr2s/vNmj8GgGG3DcTME5J+DZ1S5a6LMFRXpRHJfeF0
GQV5rkM3r80MNJhuuI+yogFGnsoCcTlVmQG+PaE4XCRtnJCb/WnVHtSWQrgIJEzgBz55c1+EiEaj
BO1mROm7KITSEMtBvFH3nIIY8j8Vy58t4pzm+bHaQIXBEogSEvAwZelS/iVKe/je9Ou4elh3SwN/
2lXX3cvN+UGB8BN8c+l5vAsY/0iC7gy1zLz+DbRv+fhgHrhI+bq5n2TODFRaIwlEUTZDX1nAUQyi
kxdiby9iMbTWL5pVQmhMEP2f330/zd4wArfHRDaKUR3V/u4wqI4SajD9K7ERVcXli3uGNTpjOpMb
JqidsdN+d/DuEc1acVDyHYx+CKbCzWYDbuxsIvS4GG757LQYGeLLXhQ8m/UixTDeXBz6hlulQzjG
7Hr3GZM+gxp9hZx1WY1IO3qV4B+eQT05KXE1SrxnzWZyy90mezE9TJUEc5d9g4AsI6p6U42zDVCb
F+60WdlhA2K03OsN2CmCwZSHl7G+ILB5xmj1paQtzUZirNli039Yk/oWH5HQTxogScnRzHpDfEWQ
2PhOJXa9n/KbXZzrMlz1e7wQKoL5pVFP2ee1qOUOeStEqmqkI3rwzXlk8sLGfLlNhT27kdviiHCx
CVAvqpCg1WBwXToHSkcmm4sPT981bmr35M+unQBrP+zE99dAzIQ02kNF0HJOLJuPSiXzYuP4ypuS
roITVF3s0/27ibhnDYbXsdr6OM7YX7NhM0sb/vKtE0VYHKuQMWM7z8JOhUwvBqBLu5mKen5sTmbE
ElMg9cHXcOzIOoSS+1PanXDH7dYzKV2DK12Y+1Anh/Jt4oKM9lvtsIHIT32fdAcKp8ZboqjEABVZ
rMFE1kGnA0mBojUvnE+gHjHQs3EjMJMGySp+Cuj0jugHGqDAM+6ZszpcIpoCyIeu+gpPlpQeb9b+
4DhG6XSy1TVzo40acMo7aQENgmsyg68PLj4rakqQ+Te8riGs+UWRRRc8SbMnDYpvglPVtTLmBsNi
mqKEHqFfCo8e7Lbu2u3Gxb3VVwOg56cXdZCQ2r3yIxWcrBBmIqYjN0l5omFCDAer1perjbP39i5g
mWY0OZpvay2QKrQIpzW+LhLfig5ZhuKYHDM00yB1eM35b3wTzoy3A/jjr8mfKM45rc20iUqanZyE
eSyzOzJd83gC9cBUYz4XbvpjDU6VHkejQegYEh3gGRPGkUK1Pj+MdJsw0rMiQ/Q4k/5BG10+h3KK
e7cqqv92sI/pJfMgTvA4M/d5G9bR4jNaAiEBdI8S8ngpkHTECG98uOpRbAijrqQylUaNTOHkIFm+
+JM/rMRT/Ngf0kVgu17EZJVCmAR8HPopb4aU/+S/HwSJTYY0llJLIzUP8Zq4np2lTJbTlzumqTJg
2+RTlXrGPSkNwUHPswBT/X3Jg/Yik5n5m+qrKj8vUbgrph4kLTcT0BgtXpSX1vgBEKuFEalZqs1Y
G9609dB3+yE5JoahWAU6JSC3owXd1eD8R7Z/zntgSxBXC1fr53cGu/rYkYRtqHMk0iViarKDghvT
5QHE8v6VVsdkaZIdKSGqvErycnEs8gptGXgOqsIeNP7auvV6gOyRrsBh28pSjsN6g6ABlzsYMeJS
hbXpVkaQWtuyw5LTdoKvvJH4En+lb9eWgk19Tn7D8usZGx6776XXsNrefNO8hlS1PJL5yB8T1VWc
l0DFNAAFDcwYwOxIkzNSG0hlgFv0qeVbdDvfOC5x7EVGGJEiV5r7FdnLE172GI4X71S6yBAL5OQW
hwLH7Pzt43ZTOrYg8egLreo2xT8ofns7+XP1sv02eZqunoRuKTb3BaK+BXtsm3Jenp55+Jz7L2Zf
ZgCoqUERDHDoEyEPG69g+IBhgsFAmDvrvK+puB1mLkpNuZZp4Sl4MuZtOWl3vkhB7A1f0gjcFy/g
c4zEBxjL4ycn1SW21ftxrC1tpHSJAk7GVwBwVYQNyVC0xUKyT/1tAphrr5oPUshcLBjlFqXHy9QL
A7dq/XXonfeNlFt9TNOxALh2DAB/dThz1uthHyPm/6/M936w16bhAJ/o/EiABMTI1UpV6siZnuQ+
rKPzHZE3GNUIcHVnC+j9xgsDQcSN7C84nrxgZBw+cnFNp3P7h5U9TorvGHQJbC5hbJynS/WmG9CM
w6FbAWPDhLxiGhkwLuFx5dtAWv1/34rEyW3SKGST8FQi1US5NUb0XyGxLY02K4rszSltJODYk1m9
xrdXR0e1v5hU/S5+2nxTqDkSRQSWNT/TiWParQ9Pe71M/phKG8GKbM2Lx4O9PkQeAcOKD5J2bp7V
+oH25cxXBwvc6bG/e8n5m7uWUmepbWho9YXJhZryFxHwvW96Ltj+otyZCZltSHqVtlCg3Hohc94s
bH1Ni+WGnmZnDuF+fTrsLSLqOvJTTmTSmK2zgiQwtdXJl5n31r9qTx3aKz3XcuvNfaNtVjVaGK8B
kcEe8xN8vUOgMgLpGtPH70CfpLfvxK2Ek/4dPcmsK2SyVzwi61oma1SUkllWqrZFNAEGuhaJV9rW
VH9n/swed4TiuJKvOgPwT7fj98DrbfvLnp8faxW4G1OAxzP1W0WuBcuQvU0ciCnube+xHxDSsJEy
QXDQbgg5SUUDkpMgyYDsMJdfloYCM/l1e23q3DVx+oly9fehPA3GDhv4nkiO7/LozyX69kmZUKaj
KA2EVqSYqgOQqakHsum/iXXNJVB8z2B+e/Y5LRmuN7qTeAusA4xKlahFHkTLRJfu3efXPB4OlvUQ
rFPOjydf7ii6+4qwT5MKnXKmvPoiah8nrAU7GmYMNcZGFUvRURggfPIRoNPRcQrMDJfQHESIc0ay
PR18KuZQmCnF+qnK3n6ekJAo+NLC9BgJJPcvAavBg6QDlOa6EdwLvj6QIfRRCgaxl56hOQev6ZNf
D6UiUBNwBgJUQjMA9eY1RMVhlpAuEiGo70N3uEvbOWNmLIZVjWLYbNrHX/OZvPm82vht/1wbYS+6
Y/OcSC+wNwfRSmPP5Q/DWIkM8tFfeBEcqM0g1xZSRU7N8h3vBuFkxVt2qc4q/4ATxeFokjdmwmAc
SHWrSX6juNy7dRMIavcZAaW3HYBsNPIV65zbWL6sK+9djU/dVfnbryzYNHex8uF2PPJxvm92zKqb
ptZG0suLoRLC3Y41t2ZUEMIrHBe4VKgLVk9Ms69EQASf9r2yG6tG4bRKDzsqR0+lkh8IP4mvvZ7e
oS+45B51thoNkeNS8qEEbsmkcQHb5RbIO8Fd1L2wl76uf0RpZdtGRjLysmY2v+h8X4dEEXteIDVC
pt+Bdas+UkT0EDCfpeiA7SZFfgtJU3NI6wBeFRFfWUGeuzEnCADwItr3GqMWtnsby0ILyDnSlMKj
UimYeAwBmqonbhELYPoQEVmH0a76fRXMD5+vbjolO8a8cIP8JqDtM9ZgWIea6CvyaqXvcr98S0y1
Vyvjg/xOdKpisPOg7lBf8AgY76a7g+mpDNXrNxr8vGBUSAcRZgxe2s+zGsOitFYPSBsFpGtd4Tup
NcaWTQeMg87nLltqCqjbdoZHGznsM6Y9Q4lromkMUozVd0zSDjUaf/ZgXjQhP5uogpOkIVsdM3L4
BIPG8vbiA7lHUQQQdxgsRbIquB0CrZ60e3z/cqXvC3L/8NpyxlQYkVUWYk2oYywJN8tf8n68Fimo
S8lRz/u6YRKXAUqrl22bCCCZSlyv14d3uxvhyfhXIAGLHf5axoqiIsa0buFXsRHJdQLpiFQ8UFCU
vj11wmIeU6Xxjqpen+qi6WTYUvsmtq1BUItfuYwYNVcDdZQ7JFUa0pYQZojGmEvqwIItZ+okjwHx
gr2J5uIYuS/+9RhIi+fBoZaxE+gwk8Ymi0se8oADBcB81+liGfvqs2EY7rIoe7ZazCuPIxeBhNnN
GA20iYr4Wv7QYDhtYDAqXFRwt8pDNZTAEHDuR+iXIjMr5EjW/mKQ4KMbhQh83DjO4qpubAG7CEcS
7r1UZtvo1NM1bFUo6P0oyEdpSTOhvqJ6UwkmGv1XLhsV5ScMAQo7JeYs4ZvIkul616NZgk45HJzY
yNkLAd6laYceRSCDEHfcckMsAxiDBjSt35oyefK/csb0WCc0+Ty2xyek6Nyv3+kAHhFPaNQ7ntUU
ZnTlgJMmm0s82R7U71Gc56Z/jKLOkdDGAA0e6uw2U3KwJEeDDchalo+g3jahDOsZsCW9NkuG4w/h
FbGScdPT8yN3s6diRXXJiPe8PVVj/z6L7x2iCpyrMoFl+hKlmfWTIDOJ2E9Zybl3K8UQ7yGgFlZd
RX8ZDOvJBBXgfFPiCVwMGWXF+ngponlciDLrdV96Loc+W+NwCWJdMAFPbXydPKWW8E5wh9YjZroi
3rtsm688UvZy+cZp4/HAdGo8Rs6S63QaTJ4eL5X8SW6fdIPDSCuxF2HVKLHEnAIGxSibZbJKBZms
z1jea1HBOq9ua6wH8ovapiBcwNLicDuFzssaKzSCHzMOY8clx3KRbTMHlKn4r3EJIIYFKArrI9Aw
WGXDwbxet2KVnDC9Bk7OrlrVNu/4meb2fWWFhgfJjaq4ZPTNwyMR+H6ROlxFZU1aDLEMpRnz7Adk
BEPMu6Zu/xLMPOb9IExKrtiewbaN8qGpq/3dRX6N2bfTYKdVjSI8eNJXPY9Q3gB6H5Gz0wb4ZFf4
BjCDBfiVDOO1zcvGDWlro92iT9UbKrF6kiuHcD6KgxpqeKQD5RWOlE1CTAb5Ymr205npJ9GtoqFB
l875XCwyC0K6SPFyzkRWEdU1cEC+wUKHAhCS62q/09R79Obol17A7QFX2ocLYKirlfSKD8RsKB24
ov7LBUHQ3Y5jIu5V8VnEIBkYJN9ZNFeQOeoOpQLBtcjGr01CvWf/FRGBAXOVgcMrAtkxUefIhQyx
U/0hn3ejcOLsxpcsVNzWSdy1/BtoujWOsXtJxbBDF0nhXbeRaU3WjzjaBMb3e2/7rf4+LB7YNkrL
pJMLYMwYriTpExyxNTABDl45Ri52VY+SGkRVdPfQRpRAWtk6XbtqjDI9QhafNdJMfjyaRRsy3KJx
eJkfNRgjQRmpJsvxZOweAamdXwPn8khAy2lJNLNe7Q7czMpRUYJm1FTrj7Cy7Al9Zknrvoh/4TSO
7mv447/xYER2wjG5CMwKqLgAaYAN9GLZ0yEVnqnOgxP+STjPc9OPUv7e1NH5UWwK2/XU2xCB4gpU
kHSoqEso0+kvoy+NHRYPQBNVE9abiFuVIUsyEvUc6ABoQBzupUQyS0Aab6j4tJEWu7i9NF7NP0fP
eN7g6kXfWEaMS5YhXhHj7LdSZd7hu9M3eTg2eKCyEsPFki0FYLvyASO9WrmX1dlKjiaMfTF8x+2w
7UtGqJdgDf+PK6IDEqTuTUrUdtGK0JNDOwFwTISphSxJ2qfv7+3s3rardkIbPvV71Kt+hZ7GRhS6
JfTqF/wdQo0iiIMgtMrefDdKCvHnjYbbTy2cGFvMBeZBI09/o+QgZf1f0dnfTELLU7oUi6GBndNJ
ITgi3+7rzRE3rXHj1RnNno7iOcXlaS33/XIT8myhY6E2IkFA9lJ4f55PE1jbo2veA8mqK1xvvEfU
cQ37CNL+/YTVlV2LPYoXI8t9uP6yYPIXfT1qeulCoiy0lIFp8+ObojBlZX/OzRFCzJSQYobT/80T
WcN5ce4JKsoJKiSxB7tkKcrk+JYiJcRlcKQndksrEGdu8uYJeKS0V4aKvX3sPUxfC2xqcpMhRq8q
Sg7vNisHwkzrSFAmMkdEXp3YvF4mFt4kia8msJwA9CoIZym03ZMesyYSvOEr7BXyd2L04K/iYkHN
RNhQZx2IDZG2xXEidwwcUgTRGiEfc71mfqYZS+k0Fxz9RcQYhLFL7iPpRvD7QTtQclNhwNMOA9L5
VkJ5Tu4QpKlr/ykYVVI0cZMqayEHrch5KIfJu3IP8HwdD09BXYAXIoFPZSYEy5HB7oGUOSWd10ak
eIt6i0uQwOhiQVa2Sta8ziXh4iqKapWBeWC03JTLoyjIONZWSexpws0hTzPYxcGOAlRO1ecxenw4
BIaTWdNwqJWxC1uU7fb3K6JwQE+xUId0ZHWYqiqJDUPobMA9H6V/+XvNso1eSugqhMpH83y+W8l+
1WxoLivgf+sVgVrqB653lQ1aEpvN6BaAAxUsWgGtc+3AgZZ4/yCC0W2vklp6YMJDcxGSG1EhKHjj
Bj/TanMiiQ2jVrnudZxZ+IdBqnqz73OyAJP+FNU7V1YT3XP+W6usqpp8MMhSV3jBU0eGvy1MUbkY
r9HTTLmuXmqIbY5mYOz7YD5XvBlXdTfAEnwD8w53178gVAN3ftmJeEgMU8M6DaOLVFdvjZuWLJze
pNNynOuUhYa334DQxwokkPBopCQv0Mbv7vFjIVYfDXhfkcGv4xefBSuK5Ecc108W4W/kW6bjd2Qy
JoN0GkPyVFTsIjKL6SdGoTE6+H4JFqfsmho5tO7KUaMCpgKmXsARs8mg0gEeo60QYc0TtgspP5id
aetgcnCRTG1JIPvcu5xSiG82kbe9xjYnbyMLpbTuDioDWqSeWvtc+xVhvRRsS/0G8yK+MursRvLP
wbupenYdPsUn8I0meWmetCZ7Mq3yf1+BuSPzPmteV1nxICm+daSWOA0OeOJdQpVhpAOargasCUHJ
mpZIZqSTGDgqUFCW7LX6vXisEcrAKRzmNrCt12WnIf6pXxo8kz2Q9e6dgoGsNDYCNYj0ftKtsPKn
rLmVMuvwEVVJWlfZ5hNeWTyx/CCtUQUKqW7YHmBj2EDH7cvRDi7EHWPpWsT8+RwooaDnsZdufG/b
/kqh8AA8yWJCdy+rMDLAnFM0+930D90KmP68xN+Pa9MbKMq/B0BZGAVKoPkBecrTe/z745VPOauM
4LM62tytEfFd8OUQ13OYpI26fUg5c2nV2tb8L5e+GRAOi/BandyuQkZV1gDYYa5FRElBrFnKJW9x
LffA2djvfZ+1ZN5EuLiTYWJ0vg9hwckvrCoPhK2EAOpqW2CkWs18R5VGmQHp6E2bXaS7KESEW+aX
E+aSdLDrdyuKGJJII0142iLqqIvOJJuOVsp8+zOr4ZJmxd8ccq0sn8b/cuiq+vPspwi3ghA7CmG5
D23s+To7ihqsiHpLH7KjNS/TVqc3r3WEAo7o4oW1LYtadjnWAsFkdy37pUcjU3Vpg6dyjjrmRi9T
avjVoW5A1x1RU+Myr2JXkPCar5eVYkBvnwz1GRHynccrtTkLX6HmPBqU4WQtdO19mHK8oaacF6TQ
VEGWWMt5R1wCj5BS3J3P2swdOXWvwvQKnchSoNEqCbknfcy3kgYtiTS5mCQTKZ6ACsXaPiJWQw1p
grB63iFmv4yU1kP8NIoSvym/aEK6mA3IWeWVCtZjyeytAdLwUG5pJhfwK5w6sFWo+LqzuN5cRUZa
JatsKuHRGbhinVDoIbyxDZzvhWVWXdZKbMt49SZ3cAa+0havNaTfkwREXr1pUCiuVze6vzZGzkSK
O9rC3RuL6x+iPSLrRPV4DHtcWYK6boAIjK1Lc0W4iARfU9cY4Wd0TWN35IcYy9AlefgIoqe2EYZz
uwMf1vHE21wGPtOdo9Q4ITfyLbxfFGSkm9VoJLDAeCUqFnN44ko1stAmC83ZLCED1U6EvKkka8cK
BaI26xmmDCbv5mbFOCIAjm5JWyrDvfeYGHhMcD98gAQ5yUIBm//y648DXUXe8bPy/SYUh0ai/4Fz
YO2ioYrFILlrp0kMZ4I8qDwXJ/ChfAA01p9vBsXMumiE+88KWWKsdAIzvyuGWWTtYcMzCFZKXp8g
R5EmmdmIPqBm9Bw7mHXHonNTQk8fWMNwFXUAUHPZatrFZ6ChRDbkbrBd44yF6Vg6lpmFjJteEoZt
BFUNMrouRn2x9LCKLyOWSORkiSdG7tjN0n6zM6NL1PpKyNmRafqWXHBJTP+n+C02OJz7nTYtfR28
yiJweOx4k+po8MsdHVv7ZDihgKmS1aR7UG+OqVsD9XLR3qKoG82WUvsZFJfnoyPI00s6cNCkA/GC
2fiIE0lJkDzpt17o0KM8p4yK8X1gRvweWTnOGFwNVCg7JycEgq7OuTl4lhSRBVxvzwcW6qXw2fZ0
PQNlSX8r9dvurRMRhMDtqtuMEBsv2x3BDp8UbXhqzNggl7AY5fkSnu1dBMIvRXCOYNfsCy7L9ihA
ii8CUnMtE0+BjeYW8wkJNU9bn+UPxbHSyGJEHhNMuUbIDfBJN2BJfNC5NaW7YDR9+k2nrSLPLhBf
tfWyAj6CtB/wd9BI78ze0wWyqUUjbT5eGOQCfFqQkOO9BUqmMBTePKulG/ucz+TllU/R77pqOK/W
NXbirBB0AlB+qouFQsNtr6xn+R0+ESMupqX+pRY9KRCx+H8vsSOEFtn4XUtld+xaDucbTj0amf7N
FBUMdxc8ieozNJc+3kTuLoc3DU2/Q9AwkMwI2pcNtDbQJwk3XZ7+32cULd5M6Xsi2JXDVRGI7L/g
/XU63a55YcwXzPjNWrykJdEKaZgaR3Ck1fDe1nDbEIxfMunCcxzJMF8imHxr1ac3IeA6+FIrx6y1
j3mVN1RXC7p+9MrMAEWkMMWCI3mZvLgOpf3f2Z4Qv512pc0UbQLX685L+t/VI9C8Umel5/s0TPOO
wOF1ZUDzu+xh/2KMopUR4xaP7lLAWjAc3kR/NALKUm+XpfpauqdDuzse7LWl/frn2P/j/S0/a7Ds
rW2fbbOnv8Jloaldj13ciLNYs6PtsCpK2eZZX18UVEFecOXTTZQKqJJYhWtPCRYHZtIT5JvTA9FU
o3aX8C6XcG9l0C+X3cM4/nigMfuxvud7wNJBl0POySc6pUxmr3+hCR5IdYdiqs1d4XOFz8AnuweT
2NFWC7kKekmzkJ5F9k7dA1Wi1RUj5yHTmoTSgKjFF6zVVSyYN9m8zxwkVFpHU0Ibvo76Gfp9LqmJ
8/55PF4ht56jOOt2OF1irp+krnVfvF91cd7BCKkq7UF2BMNGEkMAczR7nAs/j8avbgx2s7UaPwfb
lm7LIwiaoagafjmQZ9GNyj6PInUMO2r9FFqO+8WkQi7go6Tsw8MrO8QidLJSmif3Z/Asfq3oJOnT
m4tLEmJxFE3zdECrAHh08+4zXJt+SbK52OPl4Znevzxe1OypyqxFoRuKUph2Lp5+IIawFdWMkBQD
bZuQTzcLFDof6VFWoLjXuqkzY6I+xLOEZZNG5A9e+ffHqk9ks4yb96xwbdzyr1425fF0wKczskVt
kQGv4cqrAZz6MN38s54M1LdD8o+rhm34e46AfKGvLO2AWMv0+2uMVM38jY/7pGjAxRQLB1VrXrfG
4kZFA4+lxYPE9y24pnA3YYwWL0YSHKPSTXeEu6nwKfIpFxT3aDi3SXuY1x/8kOEAUqVpgaesl/Db
xKPhFSVtqDIa9oES3bDo66pOQyLWcpmhCeNeeyOOl7ib5R7c0dkeBvIazXGbDQmT4JSc6B467VkC
j/jQQj1il6GtwqwsvM4aGT6VVXLKccAwHREyuVHFjBOqwut1AllOCq6ctdlrc71S91eEVRy89SoK
+2i3+l0ljiC+x4kC9Tju5zVTqqzshQ/qcXuL/Nnu226cS9CufxhCr2mCtko1m4VxSNeZDYiGbktW
H/deB1v/7wAwuvKo0N3vtrN73yJdJHrSVj4PCmAOjoYKt/PS4kTnUmNeNHAFiN+t2Xwkfjd32rS2
yT0zDQHR1Kp5BD3/J3LYUBQowv2eq1tbYBDQV4iHZgkodUJEDmknRUcHDpOAFK5x/LRYsYsYp7Rw
OnWRsJd7bUqqhS85p2c7R0f22w2E83+l85yZD2qvSnFde2d9cCsEkdMg0OvryvN3srRkhJIJUzNf
av0kcvaMcLDfbzw64Y2hwr0LvMBWoP+/wmYAFlxf7N4AqXVvibqGt9iuk54PnLcdSwkHY9povVxF
UwvS4LcqdO+7h8ygTqNPYzO38NDb0qFTdIAv2IPRBJWvzEGDFtWti9KAOdcIPQgpMhnBK++62nGA
ZVJhCo5foLhSlYa/Za3wLtJdKh7HR37wsn5NFviqhtvS8m8R8vtYl3hb6SsOGT+naIpjbxN8qwcG
D8/TlWzogNVfwGSlDEtJwV8XyZLf45euV93pwVvgMxtyD3PGL5kNnVk9f9KwSYGkbGnSM+TzFwJx
8p7Ng5B37By7Z3Q4AyMa6rhLvDF3dj+/oLLFfegRm0WY0n7EgmYawKBBLBTR+39wikPrRUnFQJqC
nIFDvN4u/zVY28uGm4ZApNQrLvGUtcxX7lXQEg3dZbno2XGBB+Q55SEDqorqqqdlnHhX/nIRW/Fw
NAVDpAyhIu4Rx9h4isAJ9N+2TiCtzaG2r/uq7NWQ6N4qlYAcvR1SNwmJbwc8oq4h4akaY6qiLZTw
KE9tQ1tll9V2Xrl8nH0S1Vyb/jBtxIFYh1+mHQfY6X5kdRKHdgatzV6yQNfuQosPNJLa+YknGBqN
ZwXo41H0kcCLyFZxiZhUW2pPCB5rDndOYFY/T/pSQCdIaUs6ytZmF8D+lZwqkjCOR+5aT1YoYqCz
SafXd9OTFFRWUXMv+lFvNjF0nhZEzn1dsK4Hd1hmaFC+ZX+RNFa12h47VmpXd3L3pCqf4DZ7+S8l
EvGj8XHAARjAJvOSbmdN6MCp35ZCx3DoV2pGh4H6FqPhzGEkdpy6/AGyVGrlH2elN5uSCwOQMjWm
hzvtL/vsES3TASm+/M91R93XejjszprTswMa/BqZoOhpLXppbmiQWOf/j0lgeyDGDpojPsGgWtPy
CPYE0eLq5ODkVIAnvbAZT/U0Fb1N6YJQKDBWCC/urBpmI49Lwr0sDf13DfUPb4+4cTx+XT8rSWp2
0S01O4Whvyq8MPCzXi0cjCbMDLo8PYKY9CanUjCkTEuJKyCzDGwadJdnPS/KRPGSUnaUY+9waMKZ
kvfTWXC4u0WJXg/FPXPAwGh/XjbGW/Z/yeHQf+tCtSQ6Zb/EX+MIDrsv5ZE9LT9+/DNFyaSk1XIs
PRcHnFghMLzmQLbcr+9ZsY6Pu/LRjcBBo8uLS05cxpr+Maet+SUKNlDX+WtI/74pgeli/P8MyTlR
mxk62pt8LZVhKUTducaTGjBPujHsMEhpLdUpEyqsGTxZcfKVdTqixD+1nSz+3NvS04WFyjPGh6VX
1mRJaFDDYh6gzqJ1+RrLf7V27lCmt3maH2noqdOzpW7/aKmpm/TLpQ+zycPrqRKCn2m8SGauJyi4
oq19dmxHjNzmVqDKVhgT58Js9omuhQ20FBznk09HIaVopeotbyyW+ObPwfunLbpCu8f1S4X1xgYz
nBihR+mhQZerwdZxWbB6ADCAjfqfcZxi7xJ+W1BIQdzRA7RcQxlv+yM/rhvl6cpkfYobZ/ulGk98
5aH59Y3L1d1g+BvIrW7KbSwJAbopTUUd5VuoEo6g7HhOtDexo4W3IaIy83ji36sVlUoufndG+3Cq
F/wbi0XP1jGkSE5chdp+oq5907IkPB3zz34HocBTzxEwmkmycG27bm5vrvlC5nHD33+PhOXeuEKy
3sFn78hnUBTZS0B7MwvhouWOA53f07EoUhFdKkDJfhA1xb555MiDeDY4Ef19Jb+uFF7ailKlRs6X
jDEUFTEMdJtXXiEQfVgi+pe1XBzRtTMinRA8H0B7Hf/za6cSQx5b0cRkPZdWnoH7DmE7vSzqrLX2
k6FbhQiPoa0XIQpjW2ZUlVsgGDiWYi9IEf4B2z6zkVspMjiC8wcEnpO8oK0GuptnL6Hl16ZwqP2S
iivix6Mo5DzmbAvRacsuykHorNyyjbuDkgxpL8CsiFOjvv2hCXc3uPh/SwoQudJwZAxp2aoCmUjA
BnkRMiwctPH79szcX6Hs1UFRZ6g9Kr/YnR2Tq62jDzTHp1I7Gn+8MWzCSVGqgsQs50XHnC2vErCU
1vf9vEDfSVpvLrhfcUlWjwJHGL4zcv0RrBDfAFVpsGaF+IXnCXkn+ZHU1r/Wu9gSNRyHJbVWc+oH
cLUnDksrkmPs0bCF/odH26rKxzJgd2UIaRb9KuUdulBcWHmKcHet6r0INrxjnA6HlnQDwI7+jBow
aSfcJ7gu58NQgU+I79PxUSOj0PKTUj725L1y9U3rAolFMZaP5FEf/t/fbIQf2TFNPLN2xHJJRE2k
r3dESamUPrfhMI75NGJV7a32R1GUjYD7tSNy6Y4qdmtfIIMAB8epoVu8s8Y5fmzKMg16l/6jaFFi
bSuDQNxir+rgGU434KpYkqfijxPti+l8eyDGW8K+51FP+Tenar+Hqpi5kgBZ8zaNkk8NOxzazz1Q
EsaF/x47to7yqX99Yg6/DcNmy7hsxDxAq6jQYlcewyMDPqLi6CcHpcByJU3l/x3JtozUpFewz6QA
nsWLSvaS1h8JNdttJvULDNftHiLVeqs7wujT38YJyma2HckAxjy8ky8U9hDHhXBewlZtTlORRCGd
VIo3dNG11oea+rZ+eP9iArk/zp8ho055wMQmD5WaWH6vkF6/bovS31JsMsXUYEFSZn9fQPCjq81E
zEHh3XJH9253pPAmNd7BoF+zKXxhLi4sMd9uhOlQY4Z407+4BxAi/TzOOk+eopYzJeUbMl8GqoW4
RkSle43hALZWqtCBAmA5VI2jD9IgtRYx7buJwkuK62Shb6wgSetsZfJSBm1d/F93gSZtt+wzRSQi
w9Kb0jK/LbPGIxLKcEWovqdfVUghnWeHbNqqOdGwwh4bWRMj0uYNwuyRP/IjRwrFE2uBpt0iINIh
tg55BejbC46cdv58kqiWS7Dn3p+dAhbnwY3sPGwDJQKqZsUdjpoM2TGPgwU41pMLH38T2PTNiLPa
Tmb1waawCV8zdffNG5AUYwnW9za2ZTZ33wOJgxS6QOFzjX1zuSpD5z8krrXIfEqmNY2LwFYp0qQI
d1SCZvSjJ4feKOdP87bUg4deh/fAJ8IQdlKjjYrCGKlYNPKmY1RTJdJO66o3ogozItuJTDVzQo3K
HuiOB31aTuAne86I0CBe09mocKOVloPuV2zkmxxdBD1p7qvAzoISP3y2yk80/Ti51Y0HydyTgnGG
D/rIYmcs5J+8uOzzA6OPhptj6qSVBpGTQPzouxoiEl1ITuL02ky9DA4UDeYs4Nja0IyZk2fGRcq/
104NB4RWShbjf4YhRbLH5fNxkmOUexuuEiF9se6FFPWLPh5HvDn9Tp8gE/ezPftlFBCaSNSk3lGU
TKcADYl17rL0CHpi8QKmAAg6ESGvzZirnpYx0jbV5GHU+dgBGL0E/a9XVVR91yWxTvC2yIZ1tOG4
QvbZosZMJDoLkTJCt3c+C9gunHp6EPEr2DorzZv0Rx8u1zzRoMQqEoCXiOUq/wvrAziFErwpNknq
K11oBIApDLOlWwV0Y1HcufNJvb55aFaxKBVHGwwFwRl1A1UpNDALiPaNmj8Rtw2d8EluwmTQ5x3X
SfZ3G9kiRQbNinMRq7iCGR9kNXgoS5lBnC2xVhpw0i6zZfNL4+zYwK8W0OwHyzA2ym6qx5vPJltn
H9WWpoHrl/zXXnMNnopn+090nSs/YtTRAMUOGBreWPjWSOQiIshJokD2kHSCAXvWdAZSqDr2JgL7
ag+31GSVcDv+oPJUnlDWJRnGzQo+VRjVKVFXnXNzisKGToxlJ6SYU8JsxlK6Us2ZAAFXuaQx257I
+/lEDDFVX8w0Blf2rQsHjvr52XQNFrqgltdsDJgMeixcedF6o4+Tt5OLwzBmfkpwSULKaCjb2ing
3X50fX2YdDUH6FTYw1SkP5Y75g+Rbqrau18Ga/vRYXnuucZ1boUwXTOj9muRwDiQX+TdQGErtvM9
0fqknELadu476XhB4OtzytvJkF4wsYNVnb9nrECZ10j59jiiWMevmfF8WeDA1kaALNcaAj8gYirS
l1n0Es9neFXbXRT5VCAzpnlqP8DvNQNUoQouFCOzFWTC7hyTihJhxBGFBRP1m56fINArw4rTiN0H
cIT/ZyR+SJRrk0IkNn/Was/jO0OOb03ct49kY2thY6jBc7ORiDcRzhciwjzEkej7JuAK0moGCx62
O5dipXSK6YUTPA/DX1QDqvhri0ik8blEtlWjtLymEMND8exwtJj60Rxmg9egTyROz/833n/+l5Uw
JNCK5BYjaUUgv60iD9i9VW3aqnjiqFB/5j5776keedoXoc5/Cq3vDU3eOf4MKvYfTTZ/PQiOEBZf
TIhrVIZOc4SF89l8D3fS1bUAY/MhHxP26pnv+EXahE5S/Cn6nxdXBUjSy5CSOcORXUgDOJGLYuzh
KN/06Hykvb+013BHc9pWvNY15cjnUJAeCAt4LuBnPKldVTIkO2RN1D/9X5b6YrPKD0uls6h0XXG5
mR64iE5HQAB14+bQ0oK26VsX0ea9MzOksBbxav4N/Vpvk4vMb+WBtpgjCzWXMByrUFqggVGPx/zT
Cbj9CP68b2mxwoKvAWU5MNSHdigGXmf/pOCN2gZ1nEEgVBlITMXgaKzI42y63BNLBpFctMtWTW1r
6iMbcy5z9QSAqdzHJ8I9hDGfqAB/6PmJpGetSLbGt9NKkxlSbsnrGo6B88B44qC5b+NimsMXOXDY
13uOXBHDG42VIJy+ujHdLlI0PYFS2Ai1IvSWhmQzbgIev8dl3AsUSeHhrSyKTRaXb3ME5Uds1TTN
FZ+ft8OzrYe3Y7/RYpCvNIettUiFOigvgmwvaDnOq+VNwQISSdMdi5zgjc9nDwWxdfJrl4ZDvz7J
g3UjEUu1eM7apaU9hsLRrBIKFkJv/2l726pOeYjIW22ivzsxrbfQSfltBVIcz0VAWV8/AY+Pnmfy
jQMGQhlLYy3ldPfAf3hyCQDf5SZxvKEr24bcxwJ/TKkmAW45jyxyW3RD4kpnoakbpSJD/sSs4Pxy
3x6wQ1lQVe+vs9Paqzgu1YAEyQmpa0qFpkYa2lVW3M1nBKoubfZIXaDqrSaM/ggJ1fz5gLNMJSZE
PqIJbk1S97gx4IaoJtVvFskeRARJ9xH17wOuZ/MtwdVAvyC1YfhkGNjZ2mRRTgXqYfEfKiu7srY/
OTrpepv+t0AdlHkKP1G/+BkQfHbN88UU6eMbwcHj9ZdKJTPxuEWv/CC7Cf0YRF5wPdwVb1ZlSxca
fL9sO4QJHeFDk2EepK+EGia6wdZxmlxceRh4fU2MpNA2NzarXXYo8a60ZR1RKWAw9YE7p0aZa8Oa
bLasIxGbrJPBlXpcGbGGfrtdiqlenGTSdgg4RWNPsYA173krgsK3X3fLw8zTcyMRwAESRyuoaOq6
9u70PIRaYcVhZgk6dUJ8ZTnX+gijo6YR6x/2GD5tsepFiKqHsHfN8TKAxXksRUsAT/Rmgtpz17pV
C4h3uemur/E8bzsxl0MD1Jqh6xOUzylWWegEzZSh30REUSjNKfYHx5AW8j0NkyDDyG7w0OGeaiJw
RcuN9lEfKT/clcqCiWXjkjvMFfTVdRsd2tvCaJgaN5YnbRCCR5Dkvfu9D9hB3tEtIQseiMVkbDQ6
1mJM0MSxl6Pt7/o0DXqAY34qk6S3GLuCkUT3MXALAThjPJoBqa+7HD3H/78MBes/AEIriZM9QcTM
4FIAyBl5w3ZlrNocJqwGG4GU5+39Y38VtWqaLMNVdiG6RumbbWjjCvgnmKXV40ZtPE6IWavV0/fv
d1KRxwS3ilGhGTRi5g4v5+FVzNqFsztrZh4ZrOoWQy1nnZ4ncKHrNagTep+wf5HgJuaaJOxZS0lJ
ybf/2IyMJBMwB0E7Kl/vfaDSZefNVgM/tMKdWVAqH9R+nwNlJ9Z3p2W5RNodL1AX+RG0jETuF55m
fZ+RV/XvOgqKgIiUVcgn93puHZHsgWTmIpUxVgUVYyWmq1crqxGTXyT4cfrRossI1Uzs1SLbCECl
VmDwUbQGf7dvegsSO05WznGakDtSHnKNxezLjiHnpg0TWvNoGUPsAzJw4d8lVGu0t4Yd3X1hIQWF
nAACWZgvfs6H4FQ/DPMsDTD0iYWEbAemOo0IzIovZ4NQcTARubDig3LByXh7IHFtMuzDLjRyFSPc
Wbw7gwCH3blytdqvRiPTu2b7bbYTI4p3E7TWAaC2kLGEzaH3qVi2eaNmstd2tGU5L5iAGlmn5tja
ldId4pn4N3eTSm04ukD6jvFkSU0LypuFpczsiD+6IzeMov9SWV6SsmxHC0XK4cNUUwg8pj/JTCQI
CJLJ1eHFvzaFNE+4jO2eeF8gndNIXU9tqqBUzUwgjTudYhSMBq0g9NAoz1KypA0veQGZ90tTK1NX
P7y506zut5DgwDasEy6GVB/ok/O0fJJWZb97rCBN6KW0dBTs97oInq8ERvta/RPMUvWjWLDWHhZe
of+aca3B8jl7yDCaKIrrtp8tUCrlsFrbL5UZpMzf7BIS7p/lWCV4W0kc55Q3JESBk7rt29EOZmSS
b2BmxSyyUd1kVCRilVy0U6Yq5+y7NeR3Gj7Ry2z+FlwojWqRRBMgU04yRkai41IrYBtqjjkPYsy6
hVAaNK9/GzPHH/UA8VHE61nNf1s269O+PQUrJ/QlCFlfUw6d1JrPGnthOBz1zIb8jaeN5Un8P3l3
VBod7bU+AmQiGgx80Q0enetLIYC+XP51Wl7yWm8/OIEKrSsmd59HSc5VMU5zneMWwnHxOZgCf4bZ
FQoeR5wHtW4ynY3IpZENY+sWsqhhivBPmPjq6/MZ7P3ElmnuKilfC/TTbWgSfsl47B/t+Mk7ZV0v
o2Q+IRhebtcsFocfbkkCiKy3Knrc49T2gPjfZzPbQ+CyjVpVWZmicr/O1KKpiMLnzERV3b2zEykN
90NmB3Pz5CRztD6I5Dxa5L2wMZJT1l1ZPp2Dgw1OhvyWRKVk3URk5Qnc/KPzf4858Fug5UEitSfm
VT98XeFGmb73BbIgFmRp7dqJUwwY/1xKKLA051meVfus7jbDE/W0vAwvHeLHu0Xe7cvl/S8Dd6Co
D2TfCH/45iGzHtYQ6XhR3wZWhdfcBMTFhv98Dpaikt/ORTQBAnV65SS0NEKGi6T+BpOTXB7yw4hw
0XjSmysj2f/PHmo8D3ObIWeUkX88jfjJF7amBdk3skebHR8jlxH5wvDmk3x29OrFM/o2wdTtE/0Y
GfTF3WV6ybzfb3BsKBSt04LbQZeBBJUpwNhzfkdqkL43WXxynasP/FTEU9ZVcgoWsYgeiSWQJPfO
uKamattOnYsvjAYgh4I53xv6unUP8qFqyaYEtz6ZrJhGyxJ39c6e4Frmc+mhz33Ugy3X/ikBlaga
OI9FqFt59DFlFR+UGGuOOd1/G/GrDdubws2zxOYGB0efAr0FilT42aiLcO7HRCkae16f+HCjoAbN
UOYk6v8BO7bdZxTyFKEGWqgZGLU3ab2sFBuIXNItyz4/g46SiYs3/KpXakhjOU5H+FZLuAvocoxE
PjE6cShoG9zX+zqML8/HraRRO6skJyh560uWqH6oiosEWmxcFJDPjq/Y+vl3CSzzyIax7TnSN3f9
F+CgzBNtERrMzej6Na2p89UT95Ndm1YxFvNg24pZMN3X6Q5Brdmu/6wlXuJj4Vk5oZ9BYKOCGaY5
xmOuc3wV+uUqSnwqNOVCJvMgcyo3P3Rw9a0zcy7kc3Bg15ThLe48ZatI+ui6RwD01kx+XPCWz6/Y
8hPAmWeI4YrT1W/WuQOXQ/duY3DcpR5dv0MTRr3VfKgVHclyCzBk4wyvoaHFST41fDfc/sE+fWGa
voNvJBJrKa7l/EOsZUO1LRd2egDZncF41lI81OmO3bKlJCCxaiJAtrRFNiAp/gT+PdzieaJf9w9N
M3mjJQd5Ve2VJCjiTiLt26+Cf2lWTNcjx6dVIMdciheJiyOMEgaDgBkDuZaNHyY1ZWEe3RfvtPec
9kJVLEslnM2HSrNw8UM7GWg7BFvpeEYeXydlZ1YUMEYi1yDlnRpB+I8q4MEsP+1DytA+p5VnRuaP
kc4Kb7qsn+ZtKWs5k/MaXI2VQNa908nyV8ICHfgt9WX7fjl5YTmvrADxx/nF9lZVgUEpoyzrJWht
dL4Etxpd5k6+VhtG3ngQ0pIWMBhdAQgNwKKGCMeMj4DX7iWQ9wHkB0iLIS+TcCjXQzsWfIK0UmT2
JmHakF8hIFF+iTG+EnQzuQzv66ND0F/M/fNRcRESTDYYfs3GWA3O4J2PQcsbNnZRA4YCvNmXJsfM
H98xaHaISndfs2r0aYlrssEGQ2+/ZB9D9KWsaMWRL03ChxplduLk+l9hriEwn3Lh/8wHVYXDzYL+
xbeP8KlRV36lsw5qiEPcYzjwGY4yvQy0Ydqm/KfoAXJiPuqdJzKWRFMJpQRvzWGA5F5uh/WUJJYO
TVqWHaNCL50aHpzUgtBEIzMR5KWy7Cs1FkLMcxxXGYdJ1uSdfdC4YkqJYjYyN/MMcWLgS4rZb4Vb
o8iy3sz7AwVNk8vYN57zWJfp+sFUEzMo7zjh707DULiX6N6s3DqIWAjnCMv7jew6dISRbmgtCncr
pXhWgwHMX6I2cIdV6DQyWv9A+oi8KCyIoByLZs/G4iVAbIqbMgRiWctZ6yHXWYph+kUpzkFuzeTE
Ff40MRZTr1OLiq2XM1aIpcV4ajKKtmKAF8Qv//LHaGUGVB06UDtJ7MHc+N9qe/aiuP6UjcokbAkg
2h9tnSkgWRiYZVHBTJuwi1zWMi7Y2PA67B2z+wJcwCt0Sqw+i8g06W9GmtTUkbt2lBWkMBqtlhsG
9HkqeF+Osaxn2pWWkGPDNl4McCixtJka2Kz2XJBymfEOcC9cOaZDK639byV9H47PXioTFJpfcXFy
g14LZgu6uNmDaN15OJUKlgxMXj2zG3AEkIwmsU/ujFEvcLniNXE1UlH7d2elSzRNv5DeyS4Pa0Ne
9HqDHxMFoX424YJu/kKAcM5vPbRY9JqhJ/OJH5vfyjHIu964cH+C5VKCZfttKsZS39nxI0hhkban
2fEgQu6HqM6xmakLTmb47ShO+JXT3tsGfQkZd2qkQbeMEwLn/mbq5tjMrmZijXOhItGQ9hy3mVUT
JHeXIfY8JfAun7gta1psQgkGXgpt1kJDM6IzKcmVJb6rhziEZHvxnCH9A9LJr16BXSAtOuHOSnpO
OzDOYaQHnXvm27BKfxPSvAe8+42S/RpaTOYrFZ9SO5/U7o+y+zPnPWeXgPRTvSf1d6l3V3mbk+wr
R9VmZA0HI3ZYSnSNs+YAPCnw9jDMqRsMqV8xmdVZUHQxPJ5oHdLUsX2mfygxwaocPLr27Z8c8UX9
O0TFFIZoI1yCZq0NmIH7CQ78beAEw38U3HvwsOg/pqFZHBos9M7uGmBepjr+OswQmL04xt50ccCS
gJ7bi3KKg6w8V/dP05aEaQvShst1WYb2Egs5QxAmDr8w38+bm5P5jK+4qHW4K3p+8a/RRCYn4/91
3LkGgyaFuM8pemkb9faQ09q4/i/Hy6zYGTDYwAKO66A0OGeO0/q7olXOJ9MNlhmOOHcxzs3sf2fi
+lxC8eUMZbOMTG5K5YNp0lexKP1W4pVHJNCfgB57eq1ni0fmw0MX7QUb9P09yEyTl5f9k/+VMW9w
fCj4ftS3AwQKID1IDs33HvPjF7zsEKnFK8ld/nwz0xzFDpkZjp76VxBoUMfXMyLJVsVVMe23ttXf
Aa7K3hcTSWWMkf3nqMEkE2fcU9/wE3MszzfZmyznvSf2bYyOOsmRtpyCt0v0iQajFBryieh3oY+6
6nZpzq+c0KqD9XjIKxqeXow0aLHXuGp0dcXbVmcwgU4fO2l4EAczRBEexYj0mkYFFQE1i2bjIT+q
aF+Eo5KvQV3gPhaP3d6Vnq+tjyC5oHHVbqnC8irYdFdt1buePwnWSuvNQE4WIWnlRCVlZItjGmQC
B0/xaoE0SPVGkqohsKligeT5Ti+iyQrTgvL9wNSoJ+Xhc9u7yIR6/8+1nGHrsBsu65g0nEugp0P2
e0PCpr3HND/Jziup99Iq2HKB8QCZ0N/hzdIj7mK9/esPvX+8gxWGrpj3iaLHXNHvJiOP65vcil35
DW6eH0qYz2a1pL28aNdNTLSJJQZ9ST6kplfo+kjCcL8Qo52f7iwyFl70aJOLnTMX6IbaiyTF8f8C
Mvt39XQtERYdvkSq/V6oSgW1pMlZhHDIu5Ewq0he+KSivprSBoF9U7YLOgO2JklbpQfjAdSylWcz
FJEzI48ewkypqb/MfbTDyrOYmNsmkk1BfprLd6rpAYXrizq/HESqOetSzQA0KmsGVHnUZQaOUzSQ
WGqhoCCwLF4KDaOt9aO2o02o4P3clvgzrzfN88WoiY+h4Yl00UXP6h+L/ZOCWL0R+ZIRvvxe5ySk
1tx7QyFhODw7EhIVl6UqkIsmksQmUTt8JUlIcc1UTJwvajOefMBdda2WHJxM+WKw1ahErf9BXrpx
VdQ+fpGU+BBpYEouoVIHFiCba8HCwuovughr6tnWsrzTlTiWSs/HXy9uNM3dCYITb8IgHd4snxLV
Dmh7+kWxBIbg6L7538zQCn7vkYBkwjuMyszjKkYFL3pqe6Ew32jfhFufVFm1KOVAHNz6spHvHbBX
J107gf8Q44HtwDmKNWPqzeqse+URNISUC4yDH2myiFrakg/3VSfCf0LmI3JqPLLaX/yl3KuvcOea
EQcyu0/cnn5bMoRUIvIIBRF7plcnMUWXB3mTnP6WrflHkcxZYA3qIXXHOt738jrl+7FmaQJFQwpk
+BNFYxNumLNN8WiuOK/EeXRpYzt477WPYb/3aXSA/ffvBlLACWL/fGCnd/hfGLMThEPWmQUBgTsV
Ee0NMhaUZViva29wdwrbv9m7lk5x87Q6+dcGWEg926a0II3Je1PWAeayRU/bmYG1sjPb2E7kJkO6
X2pAXHoMkWDH6TScoI/dNi8ygDkwV1qx1EU0Z4WF3w1QT10xF5Mep4Ln5EQa3+n+E+IXXAcy2vfY
qmRH9alLPWbKS1G5Px8+mzdOCMNDctNzVhF+P5wC6UoGtOwshyHKnoM8z2nVJxa0DF0csBcDmJLO
3Cnpso+uz68L9yhqkt1sVHrbLGf8zmr+Bpiag64NDxhwNJwgPhDJ79M2THhaPmJ0smsCvZUm3Y2d
kREl2e/b6UOlO+SplbXHNNRm3BPxp1b8kMHNCuR308Kkjk1i5/amc6Ydn9QDYQbQR/LRkuL7vi6J
mgi4l4OT63bZtqnKPygF2DVAxVF1WJDMU3I+vjS00naDY3qbKWayjecitiLCKazgv1NOQs1vW5dw
dkHBc+RtUUMWXbzf9qrfOysGc+K3Btq5fppITgEmFtMuCmYfTRIoYe68dEuHXJlJ4EzCHMYNzwpZ
3r3hb1iqFui82YiIJso0mmAQFQGB3iBsnNXDiLLMFqQf/lEkjSiNDypMDtemx0oHAq1pbYQFNa/x
24PnRu7GopEjJ9AKIeH7eqdhnvqW/du5rX2WOxnIxfG/KnGcFyX1PwOPfKRdXjgkPMMy5TDOUqM6
JpDj47Nh0+IDk9QfxbyITT9Z68klbfpm7UPApPOoNnLJRDJBdjWcHdyRPEHyIYrhJ4lr3Wlw8vO8
Ves2rHtwXfisfKrF0Tg/6w9/6zNSF+psXpLysT1qZZI3qKoM53RCN1c2WK8nBZ4KxbRysLTi1MiQ
EwIy2grXhgdJOX8DPh0X9kZIPJalrBbXG61PtKQeBNVOMDzDjkbxOPQVXx5PuBWvLn0jEi7jLx76
gFE3vx7LAKKLhe01Jtckxkkski5gx3bTEQKtE075ZJkzHo2ajHeZZIPdVwa1ob0H3+f9XyogjaIG
lznhb0GD+6BEKnL04Jq2YJYT/XqfVg0RdBOU67te5PvZUsQ+T+bPJLMATdz5cb2LUUfcXxF/WcaU
HphmwTHnQgWXr+vbiKzjUqlVfP1GbHk7D1ycevzxTntFHRQuOsi0nUD4CsDeQDe5xGlxdvVr8mIt
q2A5hxmA0lLljWofywHkiYb/aeMV8cZvOk8CGAKFSNHHfeXhfqUr/zm2GugVvh5kI5hd7ToCAfML
B60SHPGByhwgYgbPO/46Um4gcaiys8KyUNVvw0dO7fEoCpUixbj7COlxLe7NOjCKtVyx6bRlpVah
yl7HGc30bjtmwdDxK24oOSpmK4rOoLZTF3d4uxOhpShY66K+TxXi1BLrcE9yX9xvOI/D6mfdARDV
Xo2YyApkIj0GxBelLxK36Diya6c6UESLx6c+WmuX36/RA/oHNTvOph+PDnVc0CanDuqxBRxixeT6
yXhiAG8QjHToDlRZzVJ6N3x0Mj4VKmWUm8IVPYdcqE+IeKMZhGyKxPAB4YbZiNVukvUZ4+4a0rzK
IsQZYLKt+jDIKycpT4dZCPDiPSIhhCz+go/TXZAQZZoOkn8IA7RlkzRsciDDWI8rM/Zv7TwMVzTw
gaEih0T5debrXujyGUmKk17Qm2KB2u5ddhN4JaKy4HybjjOjfTLZ5H6Fhj+9PHaZqSb3HKntucNG
pakpRzACXcAgZQHr5hTi7JH+Mtwb+M7VyRKR53oZQ1q503Iu10X0UXarTElLhpRWHMH4efyc0V83
xscnwFd+lI2bzMg8iAmabKmBlgZb1fysHcNtAuHmlh8ciukejVqGotyPJQYQE+zXCJ138nJsNkKw
DS+wSnqC4lnVPLvWiSC7MYlBH1htb/VPbrIY8g9WY3LqOL1UTElqbry1QV7LkdyXdFWEIAnmzLXQ
57BoxR74z0n2gF6Xl1yYVfqm435kWtIOGJLrju7IfYOfAJ22WcM7fMYalC7A47N30CQmOSEsPZ4O
95MbDAT2J57vfgCoinGXSOSN+fZCP6RxlR9AMAZq6c8ri/AIMt0sBT6UADQV9RBK+7gdEludbyMs
s5H1dmkfH9RrDu7NSdKqZe/QEYdw9JpiQeLo9hV+bofpGtCvqfKMBeAzbrRsX4TouC/5D/njpXHF
lIZU7hnNZP7627csSpCb/VShVgu0lPY2eL+d26f47M2HJoPSmgqPfS+AvbTHWYlUjLzRbhpAVhuM
w7tAHmMP+bSNOxgGdae+6N6LGtJPlpbh0I1o9WIGvAWBFzfdEEywAGRI4s1GonB7g8E+tuKWrhZe
4y/YhpDXBWlqFa7S11sCjaVhXkjgRZwh6fouoMlZV2AAyjRVTZV7Oce81bCTo0VYhL74f4BHxmBn
g642bHMYVHLlUaFwM70XteCC3Wy/f869acwv91z8bY5M7IPiL/fCLAOO7ix9eWW7LHVDS/ZUUCuL
zxUSUiYxJ2vPWj6n3CU+UqTpHzCfdIHY59Ml9OUfW43y+1PZUwVYKpauxDOt+87/D5vDJHILlSLU
/EXapAGFyTGRWtxlCR9yD/QLeDnZXhRUrCPUECLj/no1kqMl8FAxMt/Towaf8B+Z4j4LW+o97ZDT
HeRlcA5ej4NJJTR4zDmNnSPlGuoYJZZMIM9BeIW7NRkd49mJpJA33HUsgflyaek8Dc44kHAsGNb5
4QXmiMU0yPhdqoWPLGMwJ5IsOxwQ1TsAhXT1ILOyeTMxgm3O6s80Vx+VPey8xX952YpvDPrOXZQY
ojMYhVPSkGsCJXCT5l+zqoPO7Gqt/kdWXrl0r1HvIXZi/61nY3rolYwgZc67sU8Mgm6Zcj2rimIV
J2aJ3lTjc5wWiV4Ec9JsfD1A9r0KEo9CLMVcCbs1jTdYbO6S+dD06OBOpvwhCDG0/862dPSYkAzb
hrKwucZmGJU+exhhSTbV9UAlAKsoSbMoh1Po7+FMtlv5J6AHt4rKRr+k/Ixt6JYDA7QwL4qJ9hrE
c6zUy4pEyzbZeTU1lxcqF8gQle+Lz6XinGhKDOGD3+wRgzM3og20QeYvpmvdxL3iVApsT2qzubb+
DeXhsEbk2nu7XF3XxQ0pbJtN4umedX5Y9XPJcaRYV6O3GI0ta2tS5qmyos0Ki30icIe5ZhTeHfJY
s8snYumORQ1bakPJ0ka0UNXkk4gcGV/WVkt1RDENl0Cg2Rjo65OipC/rrpcOWB+ixnHh9evPNjTo
47Mpxe99JZTsW48qtsbCmgM0jiNf6EfH+w3e+fuwEhoVdFVc8qB4XQFOXNrmSXv6eeP43TUJoDkD
uqc7REdTTjmGd/ss2OQAyor+QCUguVyGBAWqLk6WhtGlsXAO4VOY/ZA0XAvfIF+iCozr6Bf0Dcei
UBJeZ04UBGMs/ZBZZW2LF+VXh7ktymcI1Cfppx043L2H86QDtR9b4wB/+/+/z/x9W21hED+fRZK/
0HhqR+x4usVkBhfhtUp1kr4vr1TnhygUBC4PCcnNfRVajTW3xcqTqkSpfg7gvepU0qSskBqiUAcT
zkOPB5J/fOrqeZsiZqOTx1NdyHj6xSCFAkhiYlf6+TDgNLktEBny8EKJexEKqCGaVz/4r6a8Z8na
TQhoUNOhf1F14sSMwM9FwA8MRfcJryr8Tw64IS/LZ7WiUj1DUExFM+wZeef8EbYvjAx0VHVfq4JS
+yYcVulge590cAYiSnFpWeKTpApDwUeHK77enSDKlWwrNlG3u9QW4qNkj+8vCnePbt6xfGSJ9bwe
ui/VMf67tt9XYMVOoIUgAgY9f96q1bYY5xIXTg3S8ENFtrg1RtxXtXOvkqnY/F6p7bOqIyy1N371
d1rptVMl3HqYF325xq0uAKGGmJFP7p9FdL/pS3Jfvx5GawWJOwuvXiHQeDXTZ6OvXFM8Jq2aGMuM
kSWc4WEFM0c2+k0MfO3tfaGuLrX/CdN/L32C7mtPJY7VRhWwK09Nr2CHzdf6tHzF0gMJYTRuDiKP
RCJ9388VA62/nsImBYIAqJaP5aIraGovW2svoQy+PxmheUf7sGBCfxVPa/O6dqshPtN4oqd0uIF/
jL/V4b9x0Ng+Ynu/m6j7hyrdw8Yr58c2pDYpXRR0fGSuKOfoIy0uHfw2U/H1wwpTkRO0u2zN3r/5
mMtMBPD4g6g7rVoisf3CZQr9v+zboSfUD9iA2x8E6UDyK1dOzTp3gsceysYqqrdc8C7bkqgpa0Cy
Jl15lK8i6LAfQUaEJy+npAcWSjA8iP/JlOf+Mx3N4/LMCDnh/3aOj+VjwQjZd9eh+HgQdRzviHL8
fqHUNZFpkR0h76FpT9Hcrq7gObNRnxg4xURCU4z3A7UoST2pV1THRnSsVxeY5VRryCXU4K4hZcM2
oPbEYJxKMX19VKMuQTdennpTQxn9GQDBvbeNb2CNZ2BAzmTBL7NWjtUSBac79FVv7PDZvIEt/dSp
E1S4kvYCcIjgmMiIWjLSOWc5txWehF1mmuG2iGM0E9SHbQQ8FE8EcLJnFydd5zW14YUkaGgKTHr6
C/E7hfIdovKDtsJqjplx0g3FsWT4BjplaA4l3/Yajbnai9qDyepBEpTkGRwMNGlMGTX5WxWTOs0R
1SDPzsPpBnGC+U0TqPfsNhbhTwSQX5WAp2mAo05n3Vj0JXamDl+twUEGIsfjxSq7K9kOJ766rXcl
ERaS3lI6KUfAcbGtWZ4dFVHd/079eThoM44a9u1gGkyxEvzMgC+ZX7iIianTCa7FMhDaGKszgEMY
orivRXUyb8z3CWNv15jLkkBJfPMXDjzfKx7mar/UDkzsB/MY4TY9BZcVvC2jPoWJtUwGCKMSSIXo
hIrmGWEO8DcHvXMGI/ixoDgBhddD2zKhoHIxP0wvYE+RZ1c7nfeqhj22oWs5WIKlP1bLeYVAtPiX
odyM9QpfX7X3ODgXEMxgKMeUXSsC5yEHivxMKazpsGv4XyI6TSDh8gGRFGiaTaFPTyyiXFreXWRg
zNaCjcVl7zvDR7snz9SujHQjWFhX5a9wvo3Ew1Q4DhCNMamD+jBDbvPpnVPMhqxWBzMN0q5s+/cZ
ewXJaImATVLpmCwiJ5kHaSontGjoghMIHeGmK4zEduSYwXoZanOvXDCohlJdqBr8YCMb6gInEY66
6PxxCCruZF3sb4N5g+U9poRzcycU/6iXhuq8Yi9CsPMaME5WtRZCtubW+995Y4tjS8talLVoWyeO
YKhYuvHHfPpG3l+ZkrjofjzekBTqOU38NR8cwlfayI47de1g1lmtPPC0ZaovL/XZfVv0YAyzG2gj
TjyeSgOsZ2XjNZBGPV9eBICmyso8U3YtHCEehYxE+E8q6fPHjn+i+BP7n1+4W5cA7Rm3gBQ81SbA
NbzJ+HH/d1879LY7YwsL6ScVyryb6GCwsQr9bIEK1Esox2JKWhntuinp5rfZa9YGnU3KeqKxQ6ES
cXgH8/pIIMK8cirBurgIqKA3ctEci+f140AfzcgFiOUQwam7YTI2U0m+ckISvaPxi1rbxxGpSGWA
i4/3dC0X2trXArGNpI6X+I+PCcakD1/bWMem68qewv/IaZvG9QAejybZMdz7NkU8yQ5ivEh8eCth
8tlhf2m+Ul0G/LFCQpNq/tkM6H/tT0RVd1d+Tus2V8j4DiGjrwdjR9Rc3kZbigGvEyCHHgSk62rj
hFrre+L0ahu8RSIPzH+qQCItWuzcr3uRZR/Zie/u8/wS4IdNBr5HROuDXQmcJmBSQgTQSI2OI8pk
wQqIje6A3MlJXT2Nily65ekYbIDVp0hRkqplN8HJF6xYE8S2ncskQMCOKxKvJJ13IKpfd/rhuufb
1WAXgwsqsf0jdDbIm/eSxpz+5IMiFr5rcf8S4B9Av3DYMyVpl2BU6t/SWZHDU6biEDZMIpObrsr+
DcWg3c1WdOyBLrbty6Fry9rwh89fRA2MXWgM4MhHKQuBeJ00uDPtAku7xeJt683pL/Kopd8a1sfg
LZAmt802SKtjtcgvMV/x5VFFO8/fLHolqYbbZLo+B5hbhhnfGTh0WLV4R2WSm/Lgfra7WeUYOQzj
fn5WwCZdBSi+0NbXmczxwO6jDhiSbBnxKB26ApiO1ZIATge4mjtUG6Q7c8NN1s3adLA7CJKlEtbA
m8AZ2gqLp6tN6YbeFJODLJvV4reTYVFlUkOqjmEg2RlPD3rPw/4Ob+x6K45lc6ou9hDqpA7LfMGi
veu8ZtzD9LfA3hEMtWzUt5cv5sOj69Ska3cEdpAnXQZcVRVAjQoq3ouGVG2w8Fm+633qHoqUVPto
2s0xKLQKcxLR7eK62aqX0xkM1okBdkcf+PN0UPKh+QcOQlnACFKDbGGELRPplSjg+dAOyom6VLw1
0BBKM95z8ZEaYxCouu3yQF8GVU2V8MNDDEKn4coGbyjzYVriJbjZExqQi2SB7HNUGe4SLPoytm0t
9FbDHGoskQguPkYbcW4DTI7w2ERTSVi60+rRu0evvpxrdhfEtj4ofFac9x4/rFW125txWBK3y5IQ
4ZAZ+T5NKThP3Fm4pL2oQnJwhbrYM3wKcX0K4CNrwjzliJuge7gqcNmm+fYPugVygi+7j/Z8bZ73
s97FDYyfsx7TWkuly18rpBzgWXDv6XYChh48yS/qg/sV8DzhV0822UJFDZ+JrXXzTaLA5Dmc3K3V
B9LuyigysZOWSU91hkfjvgqHn/8wROSwGqfxHJqUZOtJ8CK7Icj2t8eNFCeJhWlX0LwEi6BYYWSn
wNSHks0O/RpoPXzdkQQyXPaxYdc/nmlklk71m7rCkTr8SBraSYwujwSbwi4qFGcf2iL8mExamieK
ftQiMx/S9klhs6JBRLGU6D/cfly3QA14pWBMSs1h8sgSr2sahqMij7WNjmtNJ7LdjbF7wJF+/5jA
q6Tfs/TpVvwkuJVK6WmRIWToyWzM8HQsuVhZQaMFs+YwMTKZufpbqOBHFYIT8CHp+mjfgiJkmxtb
MLMbJN3Xvfx7X6BbFv5uIc3OaihP9+/WEcdqTyjNBkY3AKLaHCcYfQGa3vT3y6A/5mJc8oY8HxYs
Q0tELm/VHdWmXCdXCzLeii9GBlSi3fPvUILJH1a1CDmUuvxrTjVh+VsarQrPTCI8lH7xruqD/sYa
JUfaoqG3qi/6Zb3DhsymAjXxop1nNANoKU1G0RqloauFsT0DGrTzL5yP8hX3AKoSbPXZC009syl+
fdLreDx+DUanmKgVjRxx8TqIpjIMc2tP9yFOW7rfbBWLe3sPVILXaGaT46crJ2oFZ5W/GswlkYQT
/ufG5usOp2woKIX7HCk8H4P1eTe/5TK0hpvSr2iH+AKsfMs7XQ0voYHIwgd9OEdxcH0ARvtoKyka
lJIMBrAMlwJmLzzlaPABMiWuHtlqbMM1UTObNd453+Fc0buCWz3kVkcJTcB44b7yXam3rlaT+/LE
Wwg+BrzDWYuUfmip9H537DzozLSqvpJS5BoBOvSSMBQtWxaw0LgcaPWQNDB75vya3xzsFKIyopt1
tChkuevxETXWWf6WAEsuLinajhdNWXw8xSpC6My89eyvj2bHhRM90AW3V6PjBoiqOqBa5MLHHvjG
yp+TSjjkGmwlb9yxCqprhqokYqmn4fZJStznaSFu/lxb6Alc9HE3I8JBzjyrEPcAney0KPoGInll
Ale40dVvOc96kHGIqP0ov/PPVwFn5572/pXYZq1NFgqpto+MKB3H0t/n2LN9W6gG0lRK4YJsu2dk
p/t/+6LkLYpu16WVBL3Iljp7fhOuoLHj0QWPMe0gbbFInd02C7A8fZ7fqVElGoLYHenFXZeeXrWD
bhLWd6/7M8vn9cligYkNwlwFGZcfdpkkwn9SX4PRapbJivZGjAQNJsIUga31CiKUcbIus3PfoDCM
dp/N107ObTQSV/NPhmmbMvE9ESRDw6rgewjSe7Sa11EWKqvPVhb3ueBem47B7RbNCwqQQWnXse9S
0q4SYGbCTPNjUVOHlfMm2LLISC/wx37OWb9WjzL7yI3i+i4ijfRB6plaYJwIJVdnbfv+gOQacqjX
bEiZ2CaZEa00/PhxJArdQJZQFAemfVZa47JedVcchttOZjA3qusib32+ga/TyAiVdwsd5WvmdvLT
i1MRJ26EECGZFC86TOQNvZh99oDSlWYIj+F0FLJMJ+86K4GZPIsN+ukyIFtuE7EUBAkwzVGJEp7S
8GYP4RspRyyhzF9IeHgBvqdOs96BliJu9zCAsy+Z/92N3afQ9pSP3xo0hisVba5iJOt08PojzhHs
JNYSvPmuXm3mRLIw1i14pocwnvg1DtsLxoZUGLda0Xw/cRmZJg6wVJhln3rQ8Z8qdxEW1H286o5Q
B09+cnN/gw9ho8V2QmcKyNODmuf5ZbIFzcxJxm8BQuqqifHp4UY0MQyhY77cfoiygLR3jyP2/BSP
jScd9dpvZimcnj6Rz7lhD/8EK777zxzsAXPruuOaSiAt5k7uFX7H6axFMsoQRWZSJ9P3mhnQ7HsN
5PpFlrfjOEgqP33VdbKieqM/yO/9ABFBJhNcmtZkBE8LgDS16k/MfZcBbxXzZsZfGlILHJ0DAt/Z
INhxJEZkZogludAXc/iGhOM8gyur0V9Sy6j9ZoWTqYAXQBr6mQxBBiJ4NRakhlrW6rMO44SDAvAb
07rbY2Y+7WXzkmEtVG7+SRkY118DSzOpOPKvhDmQH12/I9VL9XSIyrLHfWWKsEZiDsnfmCaNxI6p
KqUHLE0jLtn/oea6kZsykvEJ1sgzqxcZbd51QCDbd4lXenWyLZdbbZ5DFPZ490YBK0hnN0tiFaUL
1uKM2EJSqHCwIYQEj2nDq9nvxuXoiFXiHWj5/fRVhds9ciduT1WM5HfLq9Z3YKFH65NIF2jSG9uQ
dWzFhiz4CAff90LsDeUQaUGDdTKlS4oNtqottmHAx9K+jd35Blre8V+Mws47MLYya8Pd8hWNgP/h
vPN1QvITuFGd0XRH3xkiMQLkGY3S+KVyZKJIhXbLUhRWY1pm31/WfdAj5DQ5eBeeFNo9kK+pgxmI
kAR8wxgsA5YU6JGlq61wM4I3Iu9x4o+K60OvaFCoTKCWlVopQi2N4eb6zSMHI3JlIfbKK883P/h+
tot7I0+Nxvb640Ix3tfvzcseq0RwRvSQEHqcsUy0iSin+JB3gl2EyClkv0SUG0eW1vuMd0M/5+xV
pIPE4kdjQjjLbkcMDOFnV1L4fj2XAz1SUWxBiggr0jUyltT1vcTsRdsMV7YKn/WYyyPcPZExCQ8d
6z4AnSjLyahuoSSCqdqbRlHVW2RI7YyEdq5acLLacaIpeS8SCMIAkJs/DGF8XWykT1Nf1Bzn4Opf
g8k+j/Tp+OTjiInxbBe5aeki+nF/bngLMhJ1x26rjk/ZADFgQ16toDrjfK/4gWjJpJzfWHwc7VrG
UtNcZWsYURjtj8DBYmx66LAzyukpOPf3AcMQuc6oX1FXXW/Qn4Ra/dv1pXQLF6Lqp+bosnCMnXMR
y2Gj4qwIIbJS0S31M/FenZiqknCMJvmw8y7cCJULFU5RyY09tfOYy3ZqcXr0TDSYpTPVX1ZZEK7m
T1nKM+JncnVQRs+y1nm6DmmEhW5FY3j8yJ/n3HXSk7NLwzeAia/uLMU1+dsLREXs1MRsGgyGDBwo
AOnzfLxFJ1Qu+/F3m0uYusceWrd6ubd/RCLV105ZPakOZrhAHTVjvPgjfn9OLVYUwyPP4krgse3s
WDGAPcpNomj/zBGaBPYLLFJ5APoMlCACQsvmDMnn9JWtKLuOBdYBjT+XjcDndLD+fjqkF2h9eHw2
kTVQ7enDjA/uPj9CfWPyQ9jfWvS4MP3z1RYJ0Qp1iNrLyqPsiQR10cWscmNliqiLSqTaX4Xzb02Q
vbjWsEtsx4vBt5DLeCbv5PJV9gZTfsZ0jLmiR17IK8ue48a3/EKr46MTxmo48r58xWZ1fHYZcMcw
fmJPfz3fiIgAO7U5LKknwgB2sNydJUAedbF1dV/PYq0UrgBnKU9gQdbTr0J66fl4P4vm4dlogUEI
VvOKZ6OVOMK0rTEONQKziaV07wFwSJxzoqZfxgNwDwdyWK+L1Ew9FEXSkKMVuy8QjeBScvLtQr8i
owO05jXsuUZEI+L9GphAvDkxQhlOvRPwpaBdcW2c8o21ckTiBDzOR70pQYGXLfK3UHZ7llNtdxaL
EGX/P7Jj4cm1sz8lnoWomwkwOPzDrn4CigR+ZO2Mbd7l/f853o3zv1yOte6C1i/DaW9E3j1kflxO
MAGJ89817f40vTmevDLZFUp3JFpIzt/Btcj7X5zxHscMer/0BEy0nDtMdge1he5TMzsr1C3XVgY2
JewQC/UIy/bbm+Nfxqowt3WvUQ0GpGWSLyVz2B5DGG3CBjNEe2gf1mjsdhKS3rqRIPt5V2Yo0MBb
ruozGxcg3ZV/e9L7tcKtx+0/TruCvWlB/wkKECigML54lEvG5iWsBn6siTiDvFsMt5L+/nca4NUP
rfXY0sIrj5XmTmEiFm3076hnmBpdQ2ycQ21J9RVLbVBQPcWe7GnTiWfb+7EngsOHAQNhu9K2UyPv
viP/2sb/K+ctjORr1Y+aIjlWaNT1GLN2vClIKoeBLBBn5osspNyFxfNQ6okQDSa+5aHqaqof+F96
i3K63zrxMxJSQ9QP0ad/CbAIXB7HLe9ANWPNk+7/Gq7FtSgX8jad9/8nILfRj3dmlcQon4Ld1Eix
HOmH426SJqFsgdzz1gl/q7T7Hp+/Yh6pNFFmIDCL/YwwZWfhKETVGti/Vij8nT1r8JsWFDYOwpeo
fqHzE7oiWjm0EuM+PHo4QEfU9/TfCOD7OsX5F6naAdkWtnJsYtXX3M8j+/NKsRNPsDXyutjl0CNT
T1tf8Gu/nkhIKi4qrsKoUGyArv+0F4symaRaeQWNE6GbY2cwQ6jtkFF/LKZSmzwJAC6OmS07YD5V
b02ERCMofnCRJLHsl2uoLOAQO1V4QACXrI/JY28Dc8q81zjcN2GIrQoUW5jeHcTN6m7CM7amtX05
Sh752cYWLFv9Xx/IkdKuRTvmKkdx1o1ZLjg3PbmGmPuFOZObGFf2PNoCyN0OmY9rjnENRYpkUuqY
qyT5qyRvtqX0EoclA4vGPTQXQF22ECgF6RabnyXR9Kzt/cFxRIhfe2exE4uXdjync/cgi6CaA785
4B14VbFCzrcv9ibTYV6UfLA3nlLTR6AAYPtGWjmSsWBtW62zlafgQZ1dY+w5NZOptB+Ghck7o1cu
xAAffhvHBGdsAWqW4boddW/LrfGRAyErLDMp6AFHq03sttkQCYM6bb9jnbLBhxIg3UwSHGajUpSb
QZ2MDmfvfu8eu00DvGAlHUrLBRI3IIUDWFQHlJjItDYdcWF7r+J6GL7WAz4uqxV9qsiapxIqjDo6
cnU2bGAv4EqGnBvbcBiewPqviHHfD3qcyradQuxQ8BPGUTadsfNIU61bIcExtNArcihQtyFYElTG
YxTh4yrSEgr/7YN6p4BqJNN7F2RqxZw7doe3OfmntzhgWHA4ENJW2sCXdj7mVjku7WKcVJMB8won
x9juxWrQlNAVaDDO0eP6wfZNhhjIHj8lTW8ZBFW0ATuBKgPFGyyFFP46FviqPOjqHS29JABiBAsB
lpoxQckda6103G8iqUGvLcdvINubrW2JhMZkgEIu6IVMSRk2j38xA77VUElxp/pNGMOTyXUzMOSO
LuM/JP7fq4cOmdprti2yzwHzpkPdAqcEgMsoGqvCu8LKF+tjSsINRoNCBN5lPDcSOL8rhax/xO9N
qDvI6hF6dvLRBek5Hgu5QToznriWHAawr+zkdx6MzvgwhsVppFGMTdsd8JE/0menq0rkMHEfEjb3
1ic8zVLDOx16omr4KfEsJMdstlUmP3ic9YqOWN2cK51Dii1/0VrGY6nDp9H+Dv66KV2Qf23HOo7m
uESpWXtNudVDU8t/AhopcjC3FXd1OdFf45pJ/elxz4+EceehdrW9UWbVmVJLhz7A6x8QONnRRI+M
tR8ey8OrohushRTntW6nreEdQJ40H/BzVvKU3w7pioY1hdDzKY2O0sZ9OrqS2XAGMeOfVD2trIYN
L2c3mo/rdYXwr2pINMA5dF8s5WibK7/RvJDTHRiFUnSVwecqDCyOK2wnAo+v8N5dl7sVz+R06GPA
ED4ZqRBdLTXIEtBdrYB7i7lI+MzMVgHejz9vTOrBdwq0SSvf16707MxZRF/WVDD0j0uneuNj2DCp
0lwPbh/eWfocqQdEGnN8W2IySsgxqRuzmAKt1tcl/2nkJ06Dx2/YjgU5nuaiGi0QtnKNrDXl71JB
QxXyeDnMqdKJup+N25gnn9GuO+hZ7FJj6cwwrliRxrY0YdrMuehzo/sFWDKHGTvQKut5b7oQ8FU6
RiV19kptwwiLItTbpGoWctWSjWD+0w5Q7IRU0sMOXbTcelmFGN9CHD4TnjxSPOMCB0XyGSR4F9Lb
e/lxrDYlNQdjD6DY5aUQybL02cIYXoWmmmytao2zawerkKL9nM6PHmt+EdBga0glD5W20ZiKnJ4A
gylADeCtRMORXlL0CUYJj805xBXmGfRWB1C9GD0c1Y8pzPxfovAGBrA1tUJMbb7wKIfwKCz20li4
Wf6QJecZzHEYHq3xVYftNtm4litF4IAIn0nT3HiYBsqChKpr7/A6+02wf8VD0r1EHNSwKDrvoGxh
7fZ9eytNrGWYWCrN5UX3MuJdYSNrlhdY2G7susRqc/Rvzy3NPzk0oXPjf61BKk/zIkJugS2n4piL
iyLIVDLgtynjlk4Hc1gOqm7kZTADnpBeG31ct3qHfJCyCWAFDBWRqgK2JhrmMSIcWl0eb5KQaoo3
gKLapMqg7QVLjB7e/C996VTnLlkdymwE1+quDK67/NeQsmKp03H2ygKZNRdZQCd0YWVE2+ZsdkoF
duTQlKB4FHgBmYrQwfgeEKF6B2Z6Ru8YCSq+/VcxI8HZCEEVUpyv74RzN3V1KFwNg9bv70pBhZEc
u+cPMO8IFz4UNHb6bmZk65tqoqPYJG91rFWlc8MQEbmG1gXoIMlEWEqfTNcJylZ2REkHir1WIPJ9
rfVPjOrQ+yy2qcUoQPvj/TmcVA9PmaZT1YTU7Lww1qvE32MvSgH1h2SGgx9zpSNG0YrRjU5QhYNT
WVDx59AeJ3ijf+Q5hXXcm+zrJh7DwNcmrVXD/Uak474/FqPjO3FowAnUTs6V/6kzpQAk08yorVjJ
Fcq2nVGCoWPqWK8cuxtoIx9XSzKQvAI3P2rLun6PJKF+nHEHsmN1/9T091MJ1EUtX6WNicSQJE+R
NsrsScrXHFpfGFbTUqR3FXTPGoTEGK9TlU/sr0+dgqdowJ7Z83f9dB2IQf0q3xtrGdzj/qsivEVb
RNnxsRg5r9UoMuE0KbW0w0KnMuZ62AzG36zFakCXOyicQr1ehu5iIjbXTJvOpCCcNfljPlcP0NKr
R72c73gbydrWjjpcGevKPCZ2nWZJBxuHB8KqIZYg6ly98rH5X2GWHwi7INfGLthHy3uUzE/Cpx9f
3rVRrQSAkmER+j/BHYya+mwn71alOedy9eFqvmKS66G11bcOe1pQjgW4b8Afzrn4mfuTUdRivYzg
5SjqADflo3yKxdVYl1sf5MAla7IK8xCd8mQpM8KZxwjp2xowBnTvYsjh2pdTqM804YAHfHj4TsRp
RjesFqQpjswpypmuL5b5iacyuwzizO5GTPZQoJML8yKIzNYBWf35pNwqq0NCG5HB2LIF5WVK5u/n
50pey9hm8iCGvVUBTIct8XkuLJTaE6RcDPZds4DslQi4QtR2aFilf3p08L4oBTufdTZjfjYanSCE
b3pxc2/Eg0gLUc+wuVfP3jk3w1ebt1oAnRixopwoUHu744mZ3rUgM0MzFjCrIVAdUgAZc4otJwKm
5nfHpHt6gCZNRHu4kCAiFx4FUeMTSyK6f7NKZWBnwXgN9y9ySYulgfMg/2KrA4oKjyq8Zz024wFg
NJlOnT8GIRp87hgGUxaKEDsU87SL9I0x4rYaxJ/ajt3LsDL8+kjvlJcsMjacdQyfXnBXKcgkkUCO
sNhWEkhL/xvKmy+xoLBBoGQN4r/pSiGy3PquG1C2+ZbuaNiIoCp3Pc8J5nGNhbr6qhKDo+X8ENv2
cohBdvx4rjC6uBQrjUsz1usmP8vV7lwl1/9t+UI6PHakg8g19asKf0vKCHWf01zpSxLA/VXRYl5J
HJlTIfY0FymWulPYTCChIaM76ivIO7BnRyITOpeUbeEta2hUQTGUMLgFLwvm/a4P3EbObRwhK1WG
/oPEmeEEda8P4wK56VkftLUpNriJ8wlJNoa+hnqsYvbZPnlIWGid7CAwa59LY5enu0yAel3VqeQR
uj980CQMOnuggVX4SsAJRUeUx9wh33VcBRaewRt7SR7g1hDV/6yX7pJQlXY+/T50qWmtikmuO47F
a6E8MnVduaoHa2GbBFDiRT6NGCUxF9UrRFQlCmoJtY3z0rwzjpNlgFi+I0LMki4+AhiZibrbsDM3
ulsfaMZViNi/2xdxiA/vBmDP+EFFEXjvrD+yS4dMTtqZDgn50xQuFcAo3R11oSty5/ZKLlhjnX6a
WvnRik9WjGlKkuIzmCg7R7D6+vV4/Sj2jgqVpkOzvaHgjUNIZqVl868X1AJ4eOzv4yIt/kuhN8gW
QVdOEOVnPNVHsgo7A8V1W/brTys+yyk2csbk+cVDHELusl44YH6hbGZedtiwexDMpYpbGBnCtdBo
LkP8o3m/LHUeYqYpwMwMpT5uEGJbuRbk/zWiFezL8ucbEBjJu1SHcx3RCj6+odk7uDfoPxwaT+7v
hQ4FnI7GXzE8F+kXvDN8YZEjEMMJnlP18jIjzYJgcSfsn1rx1ALTUma9xTdValEW5uzSQZgFRzVZ
ukYGtFbIKjavpqV9SEVIP2/kslx4zwAjIIUbbfFB/vAuQS5B7Zzx8upQHF6XsyNSJtOqLRz/beRp
2b1a3b+sFH/BXXJOY9B16NcUqVVX/GOqoc62amGedAenl6f08bAJ5vjRqGox2kvOhVuNHayJr3sC
0uHJLcXVStgZkWpcuNXyPiNzp2Euc3ynO7aZTl8fPQxJQ3w+XkTjRCC4sLFttv4WTUQjBxx24oDc
H5NEnkQu4Uzd+ASkEDjpTm73PHLlZJ0mEUmaJFqcL+W2sArz1U07DC0SFVV8zRsJbGRUV5HUIfyj
ij/Jgo7XZgoWax1Jpt8bqO3Jrc0rigaPQIR0zdtw35Ox2sF2yDWdyOZGsW56AIIToP5IKrkCU/lB
cerfnPcCxben74hRPZiW0fSolHMuScQPBfPynLE6Mt/Zmo0GqHj2jbiSqiAAtnbMj45NbMzpTfwJ
WhZX9kGSMaHeTbvs9vx8rgiuGGV4xPGurGHvEMozS8VnLXRywXk1/omIR7mMh0L1GAzxK/H11Ceg
e+7W00dNaqy9FtbXshUXZJPS/Huo+fX8iu8l1kXarc2RT9Kg1XGRljDelpiMFSFuxvV+QwF13CkE
5comxskIi+WrClhuE77KnuiEWChygGNc/axvAgxkeoQjoETNHADmXFbmjqeJnp0HTysv65cbsDCm
QZV7DD+kd3OFgbHQx3oZAJm8Z4UEY8pEOXTmemrBu6ebtUx2/qGEF52nx+czaFVX1Yy+jKxA10uP
gSoRE0AATKPYvJfG3U49jEvNVgY70wfhwiasVs7nMQM8BBHgii/Ml8R9apBpTHWqs0WZdSm+HqK8
nFwmpSegQgLW278a045fEyB9sWhSV1MvKAACY2fHhYoHH3liUzK9wJcH3NoHaizIZ29XRtZ9q4BL
P5hLjui2OXz+jWLazk/YpZ6dMxEyhrBY1ISS2wYRt3gHS4VunVLVyD/Ee4G6DWb7hVybXnyR2wDu
vXJ164IwHCqGLayYnZR/Sc6UH4y3CIPwj5HLm5y5NzEXa6wkAeetKLFYsgM5uOSmouqJR60oLPUd
Q+9ailDJiiM5fi53fm6MiRz5ixJaGvj5AP20MCLBbMVoefBh630aWaGHibuEsb8oQDVs1d3CG+/a
3eumwY/ukpPF5TJt5YEGI+zPmbimG5ATtVnlKPBWomHo8xIsWvTTPEbRym1eZp6LEqaldxsmAKau
hXB9qsvbHTETW20GYq1gp9jMRSaIucftxRUg2thCNHOnoI1oUpws312TGx2p10fbNzaK1rjNBamV
w4qx/L+N/nYFed6sR/e5uSuWYXbHjpLZW2yZLEBhGQFy90wb2jtWa5lh4qhWUZVMw7Q4zWnDOEpY
IVsdatyksXmjXGkmjpqezZzpwmtZgQTO5963jIFRAo0JrQ32vz3A0i5F934WmOumfCv6HJNlTR88
as5Lqq+zFAUKhwQRrs/MHIBVvypQOWORg2Ld5CXqo3+v2bNCfTrKcZyMRQJtD7S3iaKydpaEhIIN
YhrbJgcfFBh0Z/qrMd3Wutp1mKQZEd3LW1/6Hiin6Tb96yoi628zy1DuqdYEfbtmrRdZgdrSpP6t
VVOpV5sa4+/r6onTBKcroqWTu7SLdHwwUCvaSwKJwNdE3rE7ul41X8mgc6FAzby5rgM1XfgXnmYm
TH8TUnSwoWOqGdxNRKCAj++jGTUqE0DrIVszrF63rmWuDANcb1vwsYUrhgFg5SZvcmVz4KgdHq/R
xjtoMaRkycPEqBx1/4vkLm6omw+ro1bDjiRXNgX0wsnGg6b6A8ViOkKnoCkKmfgAg7rxgrz+epls
91l+6vJCY45qXpqAFn6lwSTooK85FnqFuE3MRLXHzkcxnBLcosFseaGSOp5BMqO/r6F7OxNip8Ep
RutkPTzWDZIdz+NX87jdEDm8ap46EgcPoKKAkm3/h78zE93A1Ks6Xb4ISC9PDi9yK1Vd4l/XczSN
aYYZGGNrdCeLLS+CdVIZAmh97cNhYEOZWYTlSBBHK711YgtgghnPysAr99vckh1jRFZ4oj0nfDvB
p883II0bt+ffsACHnRxwfh0CrRnwAEDrtMNllgvBpZJAIxDAhpbBpyuLMIlaFdzEPx1Ajo6r1Dy6
5QylBBlpwxGcQGEOulUDfehwlIf5BhJrqATQ39l2valNapDaCEz7c+sJjwHGND5BOJ4Yvu5xScMX
P2GFXqhXYG92sUR/obcm24+loZI/kwV0AxhmYon8vQPNgEi32kJ9eKqwQKuu54FzSoRN929530S0
/g7ITKpBHVWlBOvkh1QD6IYCrG0Vb13DUa7qJxrxONe0pFvGx2qftP9uQ9e0BoiK8jFYFwU/2Luk
9QaDrK3x5JzZ28ebsw/OHpE08gd0gdfc0w8WD89Ymg2Bxv9j88DhrdU9p7KPoxlxBgfGVAeKHeo6
tPDWPyfkUFQ6Iz11J44MusB1RFzxFSoWHcmGOM8c0BUu7BKID5eWXh8fDSx9m1IdixQw42j+pvmv
BcNQmSpLSTRtXfpxFhjPn/4j8eWZUG1gs1SaoE4uC0CYi+gnl0mabODlzQZpI/a4vuJGf4UkdhUo
w8oW0nOK2HRG64YUPoMKxF1qOzy1RVFh/auxbtnhBDRLjhVPI8m/nL/mK6ZAnuGGt7yG0tc1mKDA
CaXbvm5ISfaIQzphy9Nw68l93Pj0/Mfa4RyI9dcLgVAAPyJw7H7k6Gy0YS0B/Jp6MYCBtN+EdD2O
boTPw7CD/LBLWR32Jhb16SgcQgsCS5N6wKiAeN3SKhhnZZDIPjwf+7fNekb4G7awSvFfu6EyIMRR
XEKMwZIEIAsvrtXOA5Cnzt9K38LQ4M1wUuX+dh7du1n5p82i6HwfxMcrMvhnAZkH9nTYYPBBG5po
Nw75pYaXxIdYghA7+///rFMz7UnQ91xl3OXS0MLiigcZfJEcucbvCmNZ6ZN0qEVq2Q0FLnENRdji
TVMEqEx9YUcC2SZR2rSM0fq7SIiMfQoYWTEuJgftKCjaGwlMnxuBJkvX30XsNo1bJ8Ed+cVPQXZd
+MjK4vwfGoYqWrIDbnwZQq5gg4BcdEo1TPV6SOEDuCXrqySQn4qimp4/UUUq+Xyg42zQ0T6vXbyF
vRaq1TKDFCZavcm0rot3xlDW5i20XjTm09eZBxGNjg/IYWKbHW1+eyPYYFqO7wLLeW61N7zKPMy7
5wPQzE6VFDy1GE7lz/Ek1btf/00FqY7We3oUy+dubB2kvz81ioiW0NDKiMTroBUNPly6A79FJS7o
UDrW7aI8SThrRvJaHRwQaQJ/3CScMhI3XtYK7NJ1KCks8ApIzXx3iqr4+Mt0boLy1klDmOT1lADi
qV6xVYI6VGo/kFzM27Lz0dY8mRZm6D9/3O2dhv6I3yKBf0gvDJWFQ8GqELbMa2F8ICd3C79ObjaV
jMmqMGKTD2Z+5zgkirlkdBRztkz56gK1As1cUvU8XHngI3rsU08MRdZflcvNZuXNT5p+DkkFZii9
M8/m8I+MwMo+N/sVR1EzpIT5xMul+6mQkEniyyLvl+pTb3qV6DlPFJ7gW16Ho1rZVq3ugiU0wffD
dTEoRAMEsZXwwuOAIbX22M+xrCkQkDwHoU08gHkfDRCZ1/HlZrrjEidCAMFU/nFf4+k/Bbz7SdPv
1aeViU9IY29Ru4Wy4EbuYi3CiJbZILTd/ZocF0r/H+ewwEgMeDUsDyhtQz0Fz6oFeBhf4JUe0GMU
wBIJ5pjtlQCNNJkwMly67dC15AN3zKLVsuse4EbnCOtDgQKIu91o+gtDeRiuxuUw+CNk8RyadG7e
IM567axltQmrI0wxrLF5tZE1mFou4K9l0v+rwiv5K2kOfwtTiUWDybkEFni0V0QCGQ7Vs1VkVL3T
8K2NmlSkyLMxgJwyjEmRludbAuK9jBqavvwPao/wQjHR9Sqdq3zMSgJg24vkYVHJ+kjHqzbv2l84
f9eCt1wJqRZ6VnuY1Q+I+vz7OblSL1onZ67fWbcUFRvm0dtFuAYxUMAQjmGStJETO7KBW3NxwCG9
lCng9fKSIXr5NFOOC4pfpikX3KdaJE1wd4CXIsIWwi8+9TEvldn0pW5Z7lgyt+GqOezW5mj6CI8M
GCf97o1BjRJIrH2Rf5QviNnz8yHW2F56klzGrMf0zNNBD0hgKXd1EpysW8Kn3dJ+vDxUxFOWFq6N
BgPdXdGZYnVb3bhNhlzohnpeXy/JRxpDkzA6NkglJM9Pd0ZIbqOirQTrN7DnKoXVPOZjUlHvW/F1
sfPnVdxOkrmH15x8Z0gGHHsebg8fjJnerrD+3xfy+NCcvu/pE3ByrAuuKRTk/hXKlzMCI69kLZDU
dD4BGdiuhh7pxx2OF9KOwJLa3rID5NL835fxy/0qYmMqqCm3IotKh7x4griXwma1trDUPigbR4Q5
w7ZpQbAkos2JONPgSUGJmnUaNZbmpTM/O/oBvu43zzIv020ZDWxsJU0yaK6OkrtugKTKIa/1RSB3
tEw1qnuwJQKhQl82DEUWjveZVK2VL0OxDAstOjDmUT8wAgKe591UXInTJc2qW3UXpiuSGmUWTR11
ruvI84H1HUuS9ExavycP6bD2E9+ao5AJQtvzWKlMagNtXIW5oeHsjYyN6ZWwfvNBQrKJD+UOFUwa
5RltTNrwAUXj1KdrrtbYFtl2Q7E6f77qW4zSExnrE6FpUMXeA6FTJzBCXFmL+a/sy/h6HjSL8Y4I
NGkspOC1XzVOS7v06jKDyjrFSjFjOyNaohsC+YlGu95wHvBN5929wYNwWkM4ZizBIugGqVS1jG5u
HNAR6nBFk+jxwUwvnSEvqV450F8eZn2U46EMKSlk/7d+9XdnbYZ5qTsKX8EkTdYEqadlq51r9uM4
rg3s4UiIjk7F/gNESU9sbO0iaBnJgLTYxdJTDpGSkyCTEmRsBKLqR+XhoZQq0FPKdGXC7q7NDqLk
n8k7Qc2OnvA0WRBbEcTTKMpJREUoJg7MH4y5PPPa4RE9kGi46qB/sabmiWqhYmfnUs6RXajV/stR
qG0yhFhtjN2wN/cri0IVZ0BAwLJ0QOp/aSy39B2x7RLMYBzr/AcyWXJx94Y8oblgBgwARtK5EH+L
CpE76vFvAkforH4QDJBvm4L5AIZJXSguDNJSM2UPbyjPsFuNUKXhN2H/DQEQ/084y+ovs+qqL/Sx
fOPxBJr/LCUTZR5XH7Mqouj/Un1CP6Ojelsf1vgns0deJU6MpK25AOQpnTAY+xrmoOpwUnCpCvML
cOgi257cFUqHDzfH6ufwAswyJEBTgt0aZF9Ecuh3sKPCsEAkx4u6opDQDo4WerWniMYXHQ7Uem0K
uY3uGJdCYuqu1GAxVNzZwYuUR2bk4llRCKWVCGTCbOAjD5vFSjBos9XkSGgknZHw5/tdqSrIYusy
bkC1mv7CrHSr9gocfJ4KqiC87xrDQz5trntB2HyaiitS8XfrhCL2fKY5gUQIB4D5Bpj4KUZR6KXA
KHl7IEfGn4rdlBBjOELK5DftZ7Fbt9P0DBHwu4u3Fk+bMh1QX48+xVcBlWI6GExeO7cXuXUgOGy2
Eyp8ibsOkRGl89fROHTnQQG2HrfxoWoGYODiQbvY33nI7V3pOGWmRH/ITNevxs3CHMLrWatbPh6a
lgJSFvl5VrkAg33StW1OrYrd7WDLjSTBruQ5eK7UdTBl+gT/4EzQpTMS67cuYVnw97PtDneFunTb
jrrZ40UCZwWYWiLvtufn1sfH9rbCEgyq4EbJE4GYMKdTdskrmcAp/XMjMCzsf11o3MA5dYhCF8hi
cibMTAGvUUlq2N0MEjvBfboUAas0LWf/upDNqHci6pczbnhWXqAWas0GPN2TelDyiLrtMJslOHMl
FRjAKZD33DodFmLo8A2ILuE7qIMDqo3cy691t/5744yxrIKAgwIc46rpaxvPvNhjZ+pExCMjCZ0i
YRKOZ0bb/DIujGwgc+KMJDwW5zyPrR48XxVIPv9IZgvzI3bMN/i6Bq8WHRTH+cdKmwmnuZ8tnCf9
p8ANhv7L+1C6Bqz/S1gedP94cRNbkNCh4av5BaBFupIgFc44OyCpjSpovFZ9q7hIxLMsJ15VzqIm
UpRq7Toj6L3we2HKjMXQaeuyxi86EF6ykob8s2+DnV/cyyRMa4a79YlUft6zflEzX6R6el+1gFW/
Qicw10sbSkhA6R0V/vwkXM4pHga2OY1RRgwetGn8xm0MomUpG1IhLw/1OnT0cpcafs+5s6XcUlD0
HC4smghM+zUyek29vR1M7qYOGZhZ6DWyMnz2cuboa89zJ9NL7MJ9+DqjsvYSLj/JORsy7HC36d6L
uY7dvQH/ssa9GEbUfGk6gN2fAfFrV7deDlrxXSDDMwhtUWsIq+XA9meB8f+fX9P/3zfJJFVaS+7z
IhDiDYc8VducgqidfCjMNGb5vDxfaNWXEW8lNe457lXighDkxh5PuRBzFPINOLkVN80WIyGHJNpc
RTXdsOm2qpCTaKorMWSR3F8CuXPyDQQBXG7weJnpnLSSr7RUbSSGCOR+UqOgPmeaQe7I2YWPVfPj
QBE6cQj43kIGjQwkTizPC9k1VkkzinymxUp2K518E8U/hWd3W6WtJ53hFKliUit5tR/fGhdFC3h0
FLa3O506k46VTiqLtOgaxcPd2/zv8jw830lJUtV35J5i/sk0+dO5GyUOtazJJwvEJpQI65C420nK
W1Dxq9b5sLg6qViZYoNDOnt9krKOxtZHvDTVPgR1ps+dgpOvnQBdXC858zMxIZ8wSOmMUOqwrEnL
V6FPJjQxkdKEMdCbw/etiwVM8FLr3naeXMFhXGDhG4OKdn4gM7mcPKkG6qJ6S9glqaS/oaPnLKJ+
HRfeNJ5+qxJ1Fn6L3ksZTpnvgpp1CnLdln2nQOZ3PAdERZslNBFShu/Cag8BnPrKM+BG4DuZcITE
yvT5z4gUr4ysJRLWbXVV3dbT18thktpfPic/zYa5+bSAFmkYiT2JIDiVyAWpLVGFCZiczQ44Hc6v
GtH4DtPObLs1VK2QPSIK11GxW8H7ayBRR/IH/JVNfDZPVxc+HSTynTHk26ksJ7DaAEmqpLUyxWuJ
HQUne9NYu+LkmgKnUmncv7TR3aPZjX8P3A31R4PFc60BM6BoGDrHnZCPWjTP+7aEnw3204f0+mht
let+RlkPt1Q5Lk9jwrRgCrf8IADWYqCa4N8FHq3xszVQL22Sk5V1DxkVHcL/KTH4+xvFbvIhfLpX
u/h6+uNIP43kWQ8a/1qKf9V1JwxrAyyDKLPQLK3Hkv5lsoDP+MLyr4ocPWrY6exEHGCeRscjkQSb
N389+IDfR6MO8RDOZ+/2/yGwpCScX48AWnn+z+fZoch6mHR5jRPJ3ds4TA12w/V2h7HwCajKXwLQ
45uFqCCfpruroaCBJ9tPIRk9DhRnvYGXOwg88U3mLe2ze2x6hbbaSWs+otF1kbhb06n56dDVzqCD
3csBFoR2i3+gmE3rAmGI3HaZplt8Gd+Qko5CO45XYcxbIAcYxzYPIK0z1YOKui5ug8tXZ4WfkYTx
OdRqzBUe41GV3s76WNQWvpn7oqzmzL8MB7b043TyIzwOpyTcgaRR1lrX3B2qB2/Iz1rdQWdFFC9X
ewsRUSTCee0i7Se7DYRXD70ZrcAmT9yqRMt09YMS4aIqdz1NYx2HL2N7kG62jndvChSGN4oNQ0OT
c949tWiz80rzSHBXI2HXI0vLUeiRyDxlstva60nG1cjLguLxrKgfUgcYAeHo6cSZH49BBVl55MMe
7SyPNjLxvR5UkCwpVLJL2/NgleiiF6qsVCHxNQthCuzi06crO1+k4Gg3nu6BLm9af62I7kt130ss
OoKBfhjJ+hb8RaDd/XbVQ5z1z/0BNEBpKpylVWW6dZWnb5h3+7cnE4qyV+i5hh1ozfmGU4D/hGKY
ty+C6qwJQVEspR7C0isw1JBK5OIqZ7Lqvd0xltvlapleTuwwEvLTlIELblsJpXgktz8BAsct20RG
S0soYlTT5B8Qu55TJ5icPSVIbYZ3pKC7J6Da0yDACGh+Bh0xxWEQ4SV/2YLmgaVmiI+RB5RW5CKA
WEgZm31YsLrVe6Txd8BIYyeo3aKx0chrhDmPmSV3tvpQ2w+vhfCZaY3PaAkWC56P6s0GIyCbmOIt
Bhf+kl30J36zXrQ5Irf8ZQ6speylhqM8nI2JVxnAorA9tEpHQTKzIrHdEcrzFDjW9iry9MLrbZUM
+ojHuiyWZ9MD4sV041+if/Eq6BCGN4KwRuiO6PifzIlGHzslKoiGGNZkMsZ+/28nRgbJGV7nR6rn
OkhTVa1vgu+JzivckqVhbPmUNsXo4s7EBw0+QfG0hiXXnnAz/TvpOjjJDS5+SXk4K04WaFjzHVLU
aYx68MPAmnMjQHA2xRql3YiLUOilEP02dqWBaIBLZx8kiFN7OB6PJEpW2bMaps/NIgXSd7xw8xS4
MzcZJcTJ2VYiRCQ8oNDqsiE7JuynBg4IvJI4UnVmtVMBD1CHN5CA5nUYVjf55Q3YCVfjOpixAdwY
1hL76l1OshIK4w3StOOv4UdlcRRnqVa4M7GBmj23KsorgdiL0y2u47ZA4UiOS4OQu3ZJ5Lt423+v
BvKHTCz4UCxKWuSTkp0ZGia+uhEIIPgDO7hleg5c3Gpv8HVqnp9am5/Li0B9OKB4alsr3wEwhsFB
uG4tSpq/FHNgH3XkoqRlhorh+zbYRqE5gxksk4PBfhWqKeql0XyPW5CIbgz3RglfeNwKpgpGHrbM
tXOabIp2piPGNwuBRmh7vPP5V86aErPw0BpVOQZrE335SAgvnyTd1+qxrmhiQyWATxySERo3odBm
Aw0hst82rwjY/TKRzdSkc9ps5XyMQNXXd1hd7Nl2fwabOSjbhI2vojJA28GoVIzvPK1H1wjMkB5p
D9Vdx4mcaQbZUSKiPOu4rsP4xAaJpVQsAYDdE50Qb3hdQePoJaHdWfxtUrLbL4SMVa+5oXiNOwC3
e4KvC3GeoMJ1Qcc97/nbTRr7HGSSZFI04U/HhxEnLYKpj2vivYXONFW+RXgggLsTqDxErrYCo9If
VUxOD1w7OJChIov7ViW4c6DFvTPZmRf1Uq3ULk/S8JyeVhVb0dcj8tbdg9/ShoB3c1RaAQH507T7
S7Hu+5VjLT4test/wVn4orZLUI8btTcgPuifmPZKoSvoXvvs6a7uNN7v65D0fk+JU/rVoohSrcd+
+Udhka7WXY0tXUJWQp0oMvSpbUqWkRHzxgO/znRDQIrcZRBXyioxd5XRkM1tk6fIMkU9GcGh7aLT
2cc+f9dyjZvnD/1ggFTtOMPreJzscgnVDa03A/hT0yGmK8UJxlfa/CuekZLjoTN6EHh4HaIsFAG4
BLh+8ibZgEyYhBVo0PJxfdMqN/lGH7CYB/hEVLYHxBbktLks4gtXY1NYOsN9bGxS6waP1bf5Sy/E
HazelOaUMk5MFJMHYdgUvTK4OQuHuNYeSH8eN4/1OUut+fQyBGwywy/NeX3aEJSR830FwjiEn5E6
Kg0vYQ2shmZWW5Qu1jG8i9i6Ed2DH0IWofuhkWAMEIYN3hn0YaQI0lzyDMFWQghq7Eqz3Xur4dnx
DGYc5oiAdhTGsOf1HmgZNBYytTutFauqvqjIIbJqWkP8r1snnR96d01b88KtW73FQsr6tqXk/e4e
tysozTkotLL3csNN9TcUR/ys2l5x0uFpUuoJk/0lFx4pVh1YMqs+Rxp3iMvOYOkfrcABjggAKIE6
AgHs1uKu5WS2DSgX7rIVryiDPu/7YTHPto6tVln5wVi3sQzCtlJK73MKaltI1r6zw/t1bejhbhAd
7DFg22m1HRw0ZReKJOz1kiqRpWBeM3SkdQZbPj6NetwBUp7vojZRk8SnrL1LHg0T3IzJ+DRQ3Asy
cvXZiCAx5gQqAEoxwXoXfMnzwd9UktQbVhxxU1slafYLGVtIfruxwfhSbldbJ417CY/MX36D7Z7N
cOWvTurK+U2H3VHQyUaoHNt1BVc8zaK/imMnBEWtMs6kZMKW+mMtweagFyhRafeutDy08xCE0vbt
NK9AMm72a7YsEaQNofCJ+t34KH5VePSclmqiTDc5NH6chULS2yRqiYP+PZqTsmBtlDC5vNYsJy1r
Ph4dXjIf4bDC0Q4WVCdQ4dXhuJNhcFxZAzRHVKk1WxEM/ebBnVA3qHbW+pFDKB6wbkgQp5iCL3kR
R2YaC0e3tZjCydDUKDGCz9AXT7fTFd1mHC53EyTyHDU28RjCdI+0mjfCaPno0sv+Fsg9sMFaD+XW
kuO00pGkSM0037RQocxKoyZ5jH1LZDW2Oe/n5UqD+6ZX7Xc7E9tFRp69K2ioUGoTjplWgOxAlL64
xLP+Q3HLUnoAl3A3F1XyGcrWWfufAJ7Z383ann0WjAmpNZDLsq2nwd937H22G+X32u890uvAr8rV
YJWxlprCykroE2PMtL1azcONirRQ3r9UzEvSiBpWDCr0DGVTjexia8PWRYK0Xm8X2gIKTqye2BvZ
abYvHRjukF1re6H9vfJALnctuAGkIuEW6ZotIwjS6JgObHeFzzx3mRQfjaUWz+9TzJAIMQG8NOWS
DDoaLDnqu0R7zhyg0APupHRpQahQroyhC+vQi+PuVCs/w+qm/cXMmj6Z2M4F4hXSyO7Zid41BEbM
paAjuZVv6Wd8yM2X6ze/PnE1BVv4gvZi14rrpJP08atB/ULE/dUF0fvurqQONxBl7ZJneTR2RSoC
E8S5B3RLJFbjBDe3TEJaviwVH85HtmuX2N8fvjuGmqwWJdnCN+0IDuW5hHIsOZQpStHBkXSnY5go
QK8UdNZarbFPlWAfWeHF2t14MSmoHKE2SOiz3w4THVcMvDi7NfdOPzkw+vnXhGOIeBCLYjF5n6Jb
bFLptsce7H06ThJzcX6SVN5DNdXGyMOYG4jsNtbaoHtGVb4td3+yk6TOagYQ7/cadmeOMkFooOVy
vm5FG0LLKa2R+J40IsoRKqT8C1ml4pekHyBQRswNzyMU4pGN82ZeeHQuPawFlf4Gpr9kbbyBlOuX
8fHAzSRZhqxVW/g5GphyvpxyIHvrj7sO+2Hk1ESkm1BTZjKKoE1RmwG3v9HOkiq95nCBE9fgP7aK
2bkyyMjJSei0alkw+t+aXQfihrpTqwerYK/sDlqa9Z8qYRGr9v+BGA0d7IXTjLFUcSB3BN15ob63
LTMc+4nxq/ABVs53PcvFqpO5fhNTU6iVDQglKYgX0ad/CMYkfGPK74IBdGQ7T8H6GgJOea335Faq
Km+P3Ix9Jzm0P/5BoSTFiz+dzuDZhAc9fxHBjaaTec6OYux8BoQyzB4Qd2uaV+Daq4zDCUFQI2Dv
eJbPvsIKb44GoMZMdhJdbasqpi5JGS4L76p77A7WcVx6y0xWEIVAtkSHGi/JeOqjLi1g9xug7+o9
aX0Q3XuALLIkCTCOJ/72lpIXhUbn8I8SoJJlsyWPKAkTyPxttVS2IwHmAkyhk2ZaGZgw/MWiHuse
fBRu4Btdc+wI47tXCVLbm1SsZkRt/h4HW2w6pdjRgtgfPRMJ05zOc9jhTd1fHTzz9R687tJDjYSX
SQ7Ns1sfia7em2umzbAW8ZSx4okZOWyXQRlKRZlmlg+MKKLf5wDjW1nXycREmjgO84xD3zKIsw/3
WhqSNtxoRbQ1nmQkXHl7HwCf3c8nAhcRdEMw3N2dSaifjUVYbBLzjqlQzvJ/s+ZEDBogwpOJpP0J
4Fi0kPRL7cFxqeUEimQBVK9fxQ0rDOyo9MHRNIixFHyOvjnbU7JppMy1+scePfzKNX8wvgw2X71z
/DxlEy9XiSdoQQPxmNnK7mXpTP7vTL2kKBVvpbcnfthJ7vSkkh/ZPN+H65+wMNK7QbBPHku7GLTV
8lObu5OgYCA4vcpIkMdc0muTdezctbXq3/OmvMsPoNIq+Co1pfnyq2yKhFFbrECmr98xpdoaGaY9
chYVvf6yubu5MYjb7zT2SkaqirotKLtalBFQLhIju1dFTzBVgw38L9Cj6qxL5Fj9asKpJsozrs/j
outJRnpEeYVX9Mc8VYQwyMvz8javG0rxw1wdNj7XFXNQNAaXOJpGfzKDX072NtwKqa9LlPc0LJN5
hEaARlwx617f9YELAgLSg19Qy3kLIrzUz4i6eZK3NXY2EKVkd4igUgzjzuBkyWgqWosAgup30XbS
yMb5s3qnaMQbnuJY8EzpmHdevVYTRKBzke14c70gI5niL8G0QjKif2I8uoAjUS59aIHpXaIjTG+q
YrbFwwLCSJYGORsiNSWUBdHF652c85ZgxLJXHKn036P5SuuUGmTAp03mQMyh623FPCtzxsNERDSl
stOoLknFgai4z/OTp+gpcr4M2jlytQDq9V3njsEpXi0vy05Mz0E4ZN/xdlmQw/SSeJcz4dvd0LHN
V3d1zpBVozaBWH0yKTDTQJr8Qe8WXRpSEU53cVn24g8/tZmdKE5MflkTHaITPUWKnQFQ1jdsIMEo
50la24lcr4KaadsSvtN8zJ5WHHUf6uR4DeAlCa6U+CHvJBQhXh3IJOevG6gFRDTS0OSgdue+TrFN
u469mAmaKz+ZO78WHvAmTKuAiR+rpim5RPayn3zc5F2Huj3kNxz9SKAjzHhwWqkSquwLogrfxSKP
ncVv4VaMvPUjD7K4EfAbrOvAemTVXnTBBw3JNQIVNCFCmHltSKzOv24fcZPO82MuYbg6uYTgp2e3
QIzWIscjgadAJ+K9F5wdw7+SNeg05+zc1xtzs02Txkz4RjD9Cd5rjEzLu2WpchYc85eRGiC5kxUQ
sTpWArdw+xJo91mTOHnTcdfosWYthtoHryz+XO5Uisu/qqAo/lMNHefcD6WNzzVJKqPwDjUuNeWD
xeNYqOBc54N6lwgzhYkUyEup+td5TX3XRtkGO0YmNmR9FQYQ8aKsJPEN8hxQQXhnZWvvxQv3N8F6
HtF2EjoeClNpI4VXlrRDCsYolfzuJ3aNW47erxZDkVmnL/yKECNtHQGyONCGXDccz5Cg39eCdE4G
j1YTP6KSLod/tPAd5BzChP0EFwVpdhkRg3lXiDk9DWZhm1IU8lerSK/BbsT62kWXmV3K7G98yf/9
xDykU3+//Mnq6rWJjTZdof/bI/l63GB4AtUmJ0i19l4TekEOOrxDrD8gPmosqYXYWK6KVZSuR26I
eJk9S2ZmNEsYEKwVLE2hv5Wp/CzJSSfvyzpUmZTdqI8K+0uc/+bAoDOPhX+fRoS3OXv5DNyh5N26
GFk+Vl77KQEtLKF0O649JIV2/3LbGFOoRzHwjIz5fkMEShwaHAXMFN65bocERAJCwU4560GcaatD
tIJm41E4hv/oNPv+x5AhEuu+CZcUbk7YNqVQiz63RY2u/zhcHRJY/9fsVX2JGupNFgxVLN5Nd/8g
C/PAC+fy9j70H61LH2u6lR03oA6A0l75m7mLnow6qzGUevGzaChhoFnuRXx3iAx21AWcYnLMxBdX
E8/SQHNM+SCpWSHdE/vmZd3wF2pGjXmlBgiD8a6VbWD1QZHoSHMIjJsldWEBt7AkhfpQ846l+Jsv
qlCWxfNGZaIBgiYUfOovtEi3mWKmUcC7RwtYOZ3iSxPFm/gYoHg6qT0w7c7gQH+m5O2Zgi0DA6Qw
2lWka9Jg7PGExjQE5noxjdWfopFBHaVD4oWND4/Dl6a+j9p0PYDxWk/xeB305Lt4MLMWIaanmeIQ
xt5PeC9ZYOUsnVrCXw+NUDzyWfqrRyDPf9s4l48FmG4T+Bzkj+eeeXl71Ndvc8C847cNiWr5vylS
CgNQMdtrZMylSJCCyyPP2TeibK/cqijW6ctjq39SkhnBHF7XfUFOg5dwsjpSLH3mhzXjaS1CNmfC
2pdacnB/kJlE2JK9sHSeBnY1ZI3JvYeMlykFuSLicohw8SyR/cKgSji3Qo9ZH2pdOaDD76OAPN1/
0fUNM33LmjltsLkI3njwm7UI7ymA/AQXrw89LDl9N+A3d2d5zI/UaRX3e/Su0n3EV9d8tLAAZJpz
5pXjSi4DgYYSouZjbOH5FhmMRSD9arnSqeUWFZh8aXQIBRdBoROur7Zo3SvQtBp1jujCWONAhQR/
ULDStE2bKE9wcB5fKxlwqKRTSrDLwlXP9YonfoIksaZ1LoMmpgiZi+IenZ8WhYZ979l9jj0HNDJq
ouV3B9Gh6uQUbbqRq1JNSVAMa0+G9bNKboP1EVZ+/BFKj0S3R0PQ/N2slIdSf5LA3J4++odTQOMd
pUBml4NHtpBW0KeD7eD+NLOVvQvEwR4APQO0BKiek8UGDpy5KaL1vBDY6xSa4b22e31z6hU74tqv
YUEziUcZ37WGq5Zxql8RykGqnamsiDb0sc2iwxOjItKPkUxJ0pQlBXgkTIlrVlfO6XmvJ+r1yjgp
gZpqco8nQkjbM0AA5EAXf52ao7lXC9VQDsSl9LYzsc2SjVSkEvIP6hOYT8A6rna/w3NPuRbPa6DK
6qloLtZ6MuYP/7m6JHMTc4SjiiX4QxWaMC44BaPTJctxkl/743gbUMfXrziuLCcJDwBjyFP+4PR1
FFgMzlMCYJImylVW1sJWWWehHh+LzbGFrw8yXkQYgBRT0Se0qvWXu/4t7LBS2PO/vGzXiCiIq9Kx
6Wx5AIgmmvf7/wexq8RAcAmMOIcKf9NDjR3wSTUKsS9r5ChX0mfg5bw/qBG793ZI4Jr3srjQ2Rk4
vS7OaAKLcG0lDp8lS+vEJbuEm1d+bU9bGX6OeV9FXiYsYgLV6n5bHl9UUARBnkS2LN+enOsaJ9kH
J/bAevSRjwBMfoYhZeXIqcydMF8+Us1CpkVv1DcdgF7vN1dzonS93YWWu7AU3Tca4qmwQGNNgctq
L1HoVXNC13hi8iZ49XD9gt6A+hSycSi6Nxy+Dg+oZ6d88bPairRtBoaYGvKKh6IjcyMEB/+2xwk/
x7pGgH3AShKj12gRC/yb/kvfrQeKLCjxd/Fa7ee0FUCQzAYzCRvLhNytpF1R9JLYSZ422YVeT5jC
R+Wenb54svah/oRLjj3LntKK1JDbOnTWKX5PcRX3QmjUJDsYp9itB31qUtdb++wOWu5U3BTdh5Ks
hIdLNkARc6WNIYNhebJ622jPCutfYUleDssiitaITYCiTjOz/LvnbmqrJ6ohvH4bhPAqrD9c0Lon
XpnPuM4k4E9Vr/JOBi4w0kmcEAAK9/ifXbqcwiMQYpSRoS5Lh35Idgkup/t/nZQ+ffI9npNeLlXy
hXjIBasiGGRpujVk/zGRLFbPWjbEQ0XYvCJ4Ft+4/7h1VECoiZNzfZOZTz3SCJbWtSzlflAdtJqc
HEuQBDebogvAzjyl88Uvyh4/EW4tf5fqJr+/KlyJ6uOOeNaLBEYmnsmNXXg4FEig41D6R2Ue6Y9H
0oi54F2zvOXvDwj7VZPFYFP4x7agzvKI5/40zsWZ/LkZfczAi/UD7mkY1aSfIul21Uqc+y4UrVkN
mHD8pKViYhbTbajE67PhrvX70qzMvTpT0zEOKb0jdGGlSSYDQ9JycwUlZHOE9E68oxKXCRP0iFz8
LkmRrLa687n9j1IKoj4hdn7blDbIxZtSI4qnlbEgGA06F4b8ueYHHsx9asoWprPoK+pLCt8nwLC+
+zaBvJGB4n+IjoVtzy8V0ZIfr6zFDuuHP9v3zPXBLYoLpI3Ws3Z4//xjjmSEEE1qAmtF7fFD9q/d
SKHSI5t3Q6P9a3/rSYpmmIYM4oLXEp7v2SO/jE8WLH30S3GoqZxs0h3jxJrNKkTGbwNbaTo5PTSP
1wzlLawp3/tGn7veziN+UMZ0ho6ZycI8XNZn/pi6QlkwxEjCnhlf3PvVk2+JAyukVtoR6SyY52Ly
NI7KDSpyQCEy1dzakaRB2XQFEzmviOjrpsIb8G2AM3DxrEHqjfDkoiNjSJFsMWGQM6moIe2w1Luf
KNcEbQzvobRm5kOB6AO7mCaqY6GuYIlThMYa99CRJV35lPROZ4M7yhCKuEnQP1Mys5dE0Mb/3TFP
Y27/KWMSDiyq2Kmbl9XNbTYgMbmDr62NBuCViCTDX5g/CxOy7FRlSmikZHwowz60njwhcCVty3Uy
pqBke0SImSnzO/LmSOXFCLjbVYJvW2s7NShO70esZ41wV+F6itDPXAZGIJJb/x+QMbJ0SGQxJs99
EyxWATJ/cxswYWPpuc9wu6Jp65RNSA0Q+gvSHMi6MwgCLmIk75JCZ1RhyE4BgU/mKcTbGqr8EPgj
AMg8TJwF7j4rBe7ZNqtdTTYWtxogwP9aAEwFga5oP2T6kQfI6Yi6N7e8hGXf58vfP0g/WTmWN0EM
Io1EvO8kSONtkdTdNGP16LTPYTnnN5QBRY9ObGCavZ47sqcZch9A23UWwncC4g+CF1Wtav6wRGp4
yvAcDKSV3dFCQeY9O844QqiV9k2A/3SiUpiO0VwhxQ4qx7Mrhp+6Hl0dk3PChRLuOsF8Un4MU8nN
LSzYeC6hj0Z4+f+37u6/r4hBDGBRvVntkvCDcrocqEpoWo3Xv1cijNYlkfSIQiZRX7G/9Nox8TKt
xr7xzF3SEIearl6vhAsrPMUM3ORDAAHwLRo5purRvETdY//eFX1FbiceSYN9jgBQZjOJM30mqMkG
VHS8yUmYjY5nId1ufBMnGCOPiSjLkq+nnGiS5oYYSKbpdi3yFqV8Bl2uPi/bxzaVIBflygNq2tbE
6E1Fz5TCj24mvWXc9pF5NBhkOn/zb8joafkvwRE5hBG8c1L8DVVi5dbOe8/Q1Y5oCuqoF83zRAx4
0TLW9vzkUJRs182cHspodMiaemXt3eMUg7S9MfEmcAUFFLOxGrV25xnQ+J3xouOQc0G/s9Otde8T
PVblMjUyDQlAgCMlKqrootPYW1RHR+1H9IXfWgHTrvadlrY+YOXnroTkQL82x1w/p4cmlCWw8wIo
/nBCdfuvdkTMYXAzAwz2Qjlhbwqb2X1/feyb9n1N9fXjPPWEC/MG8KXr+8sNDsu/aoz5/CA/BG4q
SibNleeetzXC7Ezt+e83UJqQ1puRnEuQfwtzTFMjj8VuKf1/FEIl/DKki6TF4fejmDlh+U0Gkasv
u25I87Q+bCa6cjmMbayP60TeR+xd5NF+m74zYBp9qkO+qlhB/C3WS+pJIKjiy0o15qLiLk4YzSMj
OSTdutO8IveUi/JZ0/SZ+w+qUlp7zhVwRXHIA0j8NNAfdexnvL76PqvG0PHMjBKb6UL7KMWpX+Ur
ghmTPhn0WiAMABy0CQrVDEAgM9ZRUZ8gatr7/jdLBYMGbg4tded6PlXx5LWAu9/qf6xo9g6I9pW8
pbgTS5Lfu/FPYx1mFdqNYK6e3wr/BCeF5xe/J6bDO2568PWWl8B8vKye5lkjN4zplYwg5x4C9g+g
jcmVTtJqpanGsli7Rjbytf7GYKuGX5eyeVb8j6CZdhpNCxBrj2xIltNXPk2vma5SUhkueXhT4vdZ
MxEjidP37V0nyMJ6AxgVg/Z8KpUtWjHtDZwNXVJOqfT/l4E7riyAW9T/SwzBOmxC4XotZvh9hOjy
+UDWVwD+W1x7N2NTDWvP6rq+9PEE/1AYTi9bqWtgHt5D4TnGzcuKO2ZHtiq410JIS9aOy/T2BI+j
Y/DUg7Ac8WUuKmnzoAJoNxIMN/cxllUTFY4xrwZMtAZT0IWY2/qiB94kX5+Cdyf9/4O49uBoF07d
qaXFgkBXdVmtnt2bSrguuPxaVITZ+qkIX2dddOjB7wCBohdae/u2vtpKAaqIpgbOLaqQRCtq6aCP
IfU1xBELeVFd59Ej5/QapCxo0cFVeB4IQ9w2TMWh+HYzBnsRgS96OG4AIfyUxeB93NbbyA83Hxuo
D1TeaPgva+nAVafM6+5oOIwsSViKKLizEX59C61EsIpjBw2MYZRObh5S5M/VWZmVZ7OAcQNN8qyS
vZN1yEEr1veyxlEGq2OmatNPqvQki/qEm/+TixCUxudXXvRd6grCqotfbvkpvaGsL6IvjVPxlJRF
6YGtIQs717vSOghycmXyz0W9ybDzJCEAy08gV36q4BHlqa0dW0NeGJ381MKN4Q1lx8YR0Yx+Mq4C
/lKPk1KgifO+dLv9rPwecmhdx84S5lh0AtaEJRupN7Fl1fF0BxehxJr9k4kr6JdsmKGVSsdEiKGv
KgxpYPCWl4Wh9v6/trymD/PZliODd1pxFaHqomssGLx25n5Ph6SrCSmKmhmPJnwcy/6mZ2s90nnN
OeGPwQ7Nv7EeC8YbMQlqU1XHNXWmbkC307soj1eGhnJBGhkHM5mtj3zJXsBszDBFmIp/mOPNcBHP
atw+UHG/DgtfnVWHGEHeepo+pLYQg2RFRo/wBDvMM2DC8J59mABUj7V56KJGPb7yo/FH6TSp5IVs
7pxp+MjizOiGw67WixQ66VjDzhkVvfryYWsrWvKJbyDQ75C5BFYkl8PCJGsj33O+DNuOfqUtu3Py
gWGE95XrbUqs37U1BNgi93lI5pr7P33K+WHhyIEJgvbLkquE0e3ok8hKk3qEBIwsRVxeug+L/ro1
rd9SoMM4NR5xGorLGqZ2FrdBZ1uMalQlKoS+LF6xCuV3B3i9A2g86Mqq2Z24BdNZUFF057ZSyl/G
bkThBcONsNYQAlK5hlnYEDygZK+GYrfAuj0e02CwvmxsqtNBy01tKo1R+QaM04y5ZdNHK0v6hSeN
GjhbMra6ItzTT+sOEcP0T64/Oe6d2xoABjgQBhSz+lTAzfSj03P/NLyJNjKdrb+1i3OUeINwGEVo
GlUlP21i004hA0U35xnOJWlR50Rc60JYbe9Uk4ouYEsBg2rIVA/kU17PXtjc5BElzGwvJl0gkh/4
bG+Dg7VmcgmJbLNNfY5VE/kVJZUhe8znmlNhwpFYQ4EyA3aKevwNk4EJP3nN7M2mtyisjIwRTPeo
oNyuY4BmldbmfRhqwOsRgBpibaELNVWv0FwyjLf5Us49+EJyc3Et8ZuG+3PsT2Q+293q2TNy0ECp
dq+Q9CB7j+iddOL4ZwueUDxq8voueeMLn5HdBrxozITRkfUAkpBEnjiBLgc7euaRPR2Vv5T+TOXk
MqCfaYxG2K861jFSth6l0b4RI5pz70eSZ1jp/bOj6DKWzBjAtXj5nzRYUzdnd++6KOfcDihSihr1
iWaLHMHc/p+FSwmrqCUm8DKeQxPcvgb4Lpkb6uRnSNX60WTsxjTPgxWBUlG/lTF/GuhfwEhxyUcE
93M1gRMYcFo2yJfUJ2xrvhStcFg3SMXjahQOygQgabOH5izx50mUc/HjN7wgqMPVW/cF7/nQWfyH
HFDV1K3sQF56QxafJr8d7JGOJmgihdnVukCN3sscv5MBsU/iJSilqILYicUNfQgfH/AKPCFPAxmV
t8FaJ7x++zqgGcIw59MYKAp8UYSBpXCgIE5D/rXEJgyAezirdAQr3RM7a2fpc4WGpPu0JMHADCPu
DvVQuGW63KY/y/j4fHui1d98dMjAOgjL4541uPKetoBZG4SxZ7nOZvJgH11dclUhh7cRIanX6DnW
rcrjO7C7NjsBUNrkXDYMDQ5FMpeEQhWG9TAP5/dB63RXKF1aVfOCaJhhlS75w4PaEKt5xRJsQeJx
F2/aKCm4HzrMJI1GRxOHfF8Uq90vtk5pSyQgu5ZJN3kJ1CUIUAeMqIA6jdsEObSs+nY7UdNODa/W
oGlw+pQaW6yzoF547Tn/QclrqoQhb6O6kuZSYaDHJAJWq2fujQtBnjHCS8VrBFv6jYYFktkVRTj0
ZdJCV5TgA2BeJaR8YAj0JauSWMm2mpjCxuCA1vPbyF9SHQv21whS7QIdFdqfp3PEO1rdluwk8p/n
IBzDvLr568R2gF/mfiihCIUzUYGtoZdxH13R/Gp86NMU//pcHKGvONIkY+9jCLl+XcyozG6L3qo4
UK0kak7cOo2WIKXokNMkWrGwOa8ZKJcCBi8pby05rzz9MryII13YGBv12EY86s6pxVn8pLofnweZ
sO/FR6WyqzUoZg32BX83un+YcikD+zmPd5AMFJxq6z/xt6FBHg1vyr6i2pIWPA11/aM9wNNMTknl
irhDgXv2OBz7k+Nzi7R9NItWPqJB61OtmjwxFni+H1S2B/+wYcMevGfTwj36nJYUOgg1pkOH/J1U
9Qx7X4eCQQh8TDdaUNAIKiQRwsE4WBWavD3eMWpqp9sdMI0cF+YxAjkji7/bXq66rGw5uc+eMrGN
yieJmsk54Yl6mxcM2iwiFQHzqKJEjM71ej1ARRnX8QgfakEbANnJN8aZsLJKQjgffYQrK3vGITW3
+78b1uBQIZfF7BX5w/PzAR5Zvqo5hilEixSpfLYQUoldgjcgLfQ4YvEKbyB1ghOW+xuXmagwcce2
rIvGuA7NQLUhqOBE6kDth3VFXsP+zmJ3mIBbaxpBvBs5RlHjB9NXldRsR6/irUIbfzpeU+XCCHHL
5ulHtbBP7G2pppqbQB/74nXxgMNevh2vlykgLs7ARHZaRWHVFA7bV97j60J5dpEhTWFqwTfzvv1Z
m5a2kEnSv0+ZrZip5VK+agcpvipWxvUVgFuHntpHN3XjM3lXxxPqlW+++GruLs7hRUgn3OjT1ul2
eAdP8gcqpst0u05bAwsSBctxkjjNKmDV/NKXWXUnL73Z03bA8hxQcu3+ydjmn6xl2fLV3e8kFGkf
3x1ktOffEVaKV8tfyHlyx9mEgB4iybRp33WnUOoc98oLcUBVqBPZt9dexhDttZnYYi453srhtD1M
HcqDfUy8bLZechtuCPhftnC90pBXA02nBE6jOUCNn5auf+DAg5/AW4c5Kl6jJi3wutmEwTdgnkjH
35gBU2XHJNGlj3prfNmspjNBhGSShAxisyOhaRnOKuMR/DQ+o5uDZnKJfbF+1MJ/pftEWOXh6xcl
xKDeVRVyoYLrTnc5kOJdUBSf7ekx61wcpzBBUdrIzvIKQXpevbmeM0rTv3izu4meMAxOw+WAnC0P
NUNrAbpNA0c3Qcvfklwg0rXmoUZojlVKhHJBi16hUeX4MyiUPW9DvcjsqFTLT93WtDPmEwIPtcKJ
E5TaRMpSwnpkSnab2aM8Z7LLBWcKSo30Pxv77cayBouJX4lh7k4+tFe7QiqGT6jLoDSxClvXbhsR
lqspjlrq9jDv8b+Y5TiYSmazY/AVMe9uYaD1H7d6U7FP+smGqww+CRfY9K3A8febzN1qoxNnSzT5
y6y/OHdlwUgqjwKneGh5dXtKjLnpCuajfp9L/SM2setzrYHX1NIrgJ1U1eZvF1XfvSaoCKZxJsW6
3b06DYEgJiijdGJC7xWjfkBa5rhMKr9aTNIM8URcU1PXnaran9FJ5WjGpw3yIBQ9PNq5sy8o4ttS
n92ttWZ/A6ITdws0TXETiyZ+vdOeQHyoT0resZMsEyyyt9tDg9EP2SrHLmDGFSO4RMDVHIc/im1T
SMIjWo5yhJEmYw0uDsrVxnwhpHnBETT/5mjTL1g/QiLhlun2Qad3KQuDuX0ztM/XqioyJJDAubmU
zfAWu/5ky8+7YVK45dIB1TLa0Is0dPCcIU/oiTqncI8dNSHq/9+/dbNrR14GdZQIMRdU7Hnoymob
uwTrK29LE9CU6pzv/HKUduGF5AvjORumEJx1ZzmSOE9ttfHVr+SDm22xV2SuD3jY0cqte1daqLf0
1MsLeo3RtMpLS7MBeK6hEaAxi4ocQDd7Au5W3I835x6WLDs8g+VE1kOT+RR0kokhPfh8NqC+TR4E
GaOmV38IFCtwn9fS9qQlZ3T1ho0Qn0XpcXAHUv1ZPA7U0YYCePhM2+gN5MOTaQHxbD3XmNzHpLb0
2Ik3bZAUJ8W7mVMWHDSd3PZCZ45pWqhqYiBT34sV9doYo+1BmQVyysqfo9LCzYwvvQ7p0/zx0T7z
i2r3nsqi2krKXrxLZH2tiLYtePMQLkPAB1CaPgy9rDqnJpfvAwMb//UGIBTvro6R5CH0UuhdwTVR
LygmyA0KjdMLUGeoGlQ588WhvZso7fnxOiBQwBWSRbBjt/VuT9Qv4q8Pjdd2eGQRGDfdr+uY12Un
bOBOTFxrVoIBPg6C+2K3tesjJFSRUKlG8Tox2hswjJ4PX/pnLLFpfgGmxPPfFkrKiXlVgp0vILY1
47BPqLKZ3TOVdj6qbAwfK1E2Rt5aI3zqE3KJ4vr8LpnM+EkV6yXG4i7JPmf6zS65LJJ0qe5Edv6e
CbW5Aghr6yXFlVufHaJVBcm4S2yNCfkgSyU980owm7Zsm3mBHWU4gNjyo2QsgrU3Ufey9K0Iet84
XUoVv3cBo3dS+viJwTLSUPiNZWrcGE22lhZvF+ZAJg4rvQ/mBCUwbtZ+12J1+oIXctB/LqLEpltg
qgU8tqXyHTXV6RyIsBtR/jI+gusbvmSujU4zmPJYHaF3+Cs37ulNHzaQjd8FAhnnBhjnw3ZEevB1
RUeIfVaqsHMD8lqJQ2wYTNdAws1584qPZIAFSOiBr4HG81rLRrVFKzi+u4L9tK1+pW56jsROAgQL
A83M793wG8O0X2LDZaoV3kFqI8fwxYG+kdn6LiKrVXgfJsZ7kraZ7x+IJ33a3DWPSnA291dhVyLZ
ySohjMXunookDDwZZcnIf77l+xCc1qCOc4Knb33iAdhG7q6+dXQ1ZPxepLQ/8XiVfP9HoPQmTEin
4hhYaXJF/GvifNnzsH9yDw+wqDsma4uJ0v6C/HTjva/Lzvvmp52UC0M4NO4MuLCS3sg2gccQqU3o
FQ76INScY+YX8v9ZeRSETEPe2hnrmxLVpCf0pfF2/0rGjtoHoYHJzP6W3xqXnPg4RxnFPruXVWyh
XFu33LUfdP+2EITJs3yU5rc6pvO2gU0riM4KAtYBkvEyjA+KdT7w1dqqC0lO6IjyTOH+Wi1nkRQd
XUuaTNFgRvveY3cZANQpiXkUQybcN20Uunuy9/PF3oeh12XOd4SEaHIshk79ziqnRCif1JMVx9Do
0gy9ulkyRtl7PYvJaM1fnAHfhGzrSjO6yXauL827Bo1M0FPx5t6SByMvLeZg3g4bNMK6hmIfoG9l
AAlX0jxlHHkbuSGtg86nrl8hVgchJHGcql7pKAispI/KIU40vt6LfdbzpUKh+ojsoytEz7MvD4fF
yGTCVWl8ygs5we5+ACN/ERFrT6udjMt0KeQFAyox+QSHHpfIOQoX8PprMgR6mRBTFs2VCHQ0dFPm
VbdOkXZaGJueWZXBNKs6dUC2iheKMX9dwM6Ni7Dk7fNEkVfEHNwaw+lVVcCPKhu+49S9gxI6Dggv
WJ6a1jfqOTTcybWAOD6dteeZ1NYc8VojL0BSBqNvx89HUj/l8rvyq4dNDcCwQt8QnQ9P2q1D8ocj
21ST9PUsoUhxlD7RGhRB1O72ychPimfN5EHTOidN/ADTYKfmRKscfSVTBjx0T3wtFzDP6hBnvJZX
s34dIWKy04u8vvoLtJT1q9wg9yyUTocsFRfh+EbX41ZD/19IytmagE8fWUKNj1l6UbnzjZq5gRui
L8X4NFdXKqmLFdQGElm5D9R0XoUgoeft7RG9x1Lg1UlEB3lb/bXalisW52bpnrqDDFg8fVnIW0pt
r9cpRSkq+0RF0ZuOCwrxezTICvTcYlzVEuMqIA0otmt2+iJ3z4JerUIZfS9YCrQOPAdG81K29MDa
4C+mWwlngTWdz07iyl6t5UNNj4KmFo9S54qJA6BKYAfyHXV1Rz0YV+37AOQJlc/oOv99kn8jCP3H
I1J+8i/c6+s9YPJzW3dUyDDw5MVawI6rGr+GLsPJjJqguJKzaT7cyJKXG7bmWEqxaLKRnFtxP34t
2BfKvhl7AQ5lXKGEnaqdvzy2gzSpqmJunAtWr6EkBcaWuDVA8akuAf5s0VD09+nk71ociB0pbA1/
FarOopqMFhkXna+ulXW1tycjQlxSQ5pGxRcrnM1e2Ls0grxwVzT58gBkuP2jJ7Zj4A1OUPDckuGJ
APsYuSfOiyU72sfq9sRrVZgG4viC61qmTBm9lSnPglLcdEWz6MwvLY+OYRjdeqA+iCnLKXGh0ZSG
04G6hrEc3oHB4y/QFSrtKPXhSspqJ0Bro+HL3779eiHJ1uJtf2c75bKJpTIASk1/y+P9jRZC+MgL
v/rXvIBY9RoumstqLWv1hoWJ/1Ckb9E/gjvZ1bHLmfWsug7ybnEwWhZji5m4ug4kNkqSdqimTvoF
PJvEeLVCzY1guEd9qh5OCDOgfUiscuAFEvUjkpnrSmJK6ByMNDEZiYfHBZK/6nfqgF69PFB4eBnW
nzwanKAP688/cflIpCM5TMdFSUabU/qw9w2La5gWtbdD5fi3h+t2yUuHEG+0P9CU9DPdtfTtO30C
cM2uHa48Uwd7JqJXs+nfBsLSdUZ7K5x1B8qjQR1tlXext8nD+/7YqzYczTgDB70xmP7WzqgCDnqw
g+/2Ura75xUbvM+1yKT7vkmcJ1JMRyl7UOR/JOjWNVmNsRkAhfViEBCF2V9yUMwfUnP3lRkbAvZr
3mZrj/SDfq46VzxwrXu9enxMUA36uyruuNVrGGZNyPjuzoQ8o9u3IyHnHHRfJxZCUtwFFNBV4XKo
KUX8l12Va/STuwA5IVo/uZiVyMzpqHe9mgIcL8YvS0aQFUfX8EjPNqSxsDDV9CxS3mkUFTVHSsQ7
1XTUbU6VqWfn/ZPS2aMmEba2nwteba1MxI+B0kt8Oso2HM3pmUMD+q2nsv9bDJ5cQ3VVDYtD2VrZ
TSM7g6av3bmBbZIGhub8RPicS4CyXzGeIDpsLME3u8veleERc8tOwdhp1Fj3ST8qASXIRvVTxVpH
2R/Bi+NqJ+5nk8bEYu4+1dCHb/J+GWU0UvtwHUXQdzyQivVSkQARGA4GttFEEsv+tHf3x0HmyLMX
ZQqqyZxc3gFHKsrfceh75PqD+uADbLshaajpCCDMI5FLPqEmjsDRph5I+1fZmNfQXiraVfuZmytI
UQ22+Gx3GuBkUIC2+oGV+U6+mbbYOg7mbJuVVh2d1l6Y6yqomzRkYGYylYVZ1xGXNnqfku1LyREG
SZpLlVr2q6T2LPFaUffcPHh/D2dTpBwUlvF4RhP/9lCH/DsZ4zgdcpkjYeSsZPuQmR1rvkzfY0xt
zalVtg0i5an49y8e3XvxNNbtue40t2Ussz/UpxlRnEkqzZvANWDgvPACPnIzp+6OYLY0ns84/jLx
3ym7SOhVYRS7Pfgb6ixMHJkvM6HZI56utrM/nEpc1p/sUR0iITxOUT6VRNHzIOIdUJmDQ6f1gUxx
NS1PRPxSpHwLtH23gqsFrDfKH4lkFQ4zLVdAiQJyrHj0e6O0pFWOVWQS2l5whCsGY9IkqjMrKdzJ
2rJAaFX1PHtAC37sL5ud6CZnGnapflUTvA8os4jhUb2R/L4JIXUWaBIniK9HgNErH2gZYtJs6LPw
JHMUxv7AQ/IgCS2HhWaBCG2TZNcsw1Rlmy2N9uBCwVQKPQ8XyxIRsXLaDlfmm61npNgCVYw5aAbF
ottT3U9JBH+y7mtaDGXW+73lq9Zp9zdm3iBp3hzJ+x4c2No/omB6imz41VOAbCle6iibjGohBgYi
XOJoNU9kHCGwmvuR+4GS64W00WQrBZaNJRPw+JFcAL6jPPcU4rY2Wf0kBU2/R2DeTFvHeuPl2akl
pnLfQQpYI1wcA+T+0QAkW1H06KNcEgUyIT80EdgTaK0wD1YRwrMALMEOtqW5OIQqV2vG5KMnHShi
g9y1XvL/XxiGK73IIRTGBPfqV+lQNvJ1BkLngu68MrkN640+Mjq4dagidRWdEd/acR4RilBRSSOd
kZX8SWnWJZw6TTKhayJFBR5/uK5+WwuJLM/3+x+UHVyGg6YPR/0mTgLBNDLnmPia+KFDDRJZtazO
hfWSgGivWtRGsRhHg/MaAiUO3fSJzXS+9tCnD0diqMueFSg04MjbBRK0CwDyDGaWtu1q3+oOA2jP
AECHVkdxdal7yofq52m0qKNbMgEucHksIC2yo4hdM6GEjsuTVd8ya8jQkSR3BnKXuBJ6OlM0S2tP
nIAVkOMHjZLVN55LYonovJKOyEycHVgoGlAqFQwdl/ND322Leg+yv33F87MZfvVVEmKOGx8JMK1F
n45EmNDerk5wkcrsJWYCvoImhT0Ne5X9SZpI9H5qSPIklciYZqSiAp76jSLzXihPK1fARTtNXp4s
QRcPtosnULK1RQRQrYogZAQvvp5GLg8irWCnv7RZ4Vf9CDglAK1l+Y2mIZhJA94D7aRHaXQ6P09Z
JF/xrHLWoLag8Y3l83bPg64PBu6G/R3iNPaRIYb3OQadDDEF6GRsqeP7uwLmsFrY6TmFYZkwXdKX
mo6aSZ8my5lHz5C1267z0T0sekCTRspHGr4kHifyYprWAFKRixKkyBsKwbQu4gG8MBU9coi4Zi/G
DsHjzSk4sZaFrC6PLZYUL+C7KERwBxnVI4zXzc6Lq7w5ufI4t5Ev87f46CYlyH/MxfQ0fxd4h2+D
7m69dFmiNs0Mmz7WPD01//p9C8HEnqTEXJbpz7GHhh0znyQiHz1Xb//wdlQAalgeRZXNTaTjtF6M
vfUkwwOusAuEzb7endF6WP8J349schuQUkRNbF+Euo0qo2JYkJL8akrzUBZIc28H3IfQwJXG1J6E
T1ZJ71bzfZMILal/qGZXIdhAwSKR9N+kNlq9RCb7usZfTK9mmIxHkv8INIg1eJjF7L7hqJB7bel3
Z2pf86cwXF++o50G3h6hRE8Lv9AZH2s3zpLsavBLa2yy77/2App3Hs3b6FJPBvaKCfCltszx29fr
1IkCLbqarlsECkrsejLl/NFZrxpppqIgrndJTymWxj0Puxs/+gvuxOdppHGDCli4H7B+85aeVyjO
8B6tTMWcLu+NswmqRGq6fg3jFLBmyG+xlIp+6N4n1JGDApsj7Vp/Kmve++EAWrku3W+5eWyfaXr1
ITbArxRLihfaAzboTOnsPHKv46Rz6eeMHohIMBWIA5uIktHlcyOIfJOCMIe9UcxIdTnXFkpXnBwE
YWp5rCU4JVDhPVoDAi4xgZoEi8TZXDIy9Pi8HBkcev2phTRaggSkxj/82x4+BlHJ8D9PP8y9sm4z
GA6iotvEnRMWj2SlDfgyEBQrq6LDot8uue5DWrW+fXUJTPrk3Q54wbWnMG/N02L49s8e7PhRRC+/
mfVmoY415/6PrYADqBMDPHxmSSooBY9ngI3cuQ0Q8MkfYPZHcY8TNCuGSX6RcdIz9uD6XOL88iBl
evLpPi6C4PHGnyzBQYqiUgWO0HXZw76bNimhXxVSNL8dr4YsFnTPTPlGriuy0hgu57HzOX3sfYjv
gDoY7rwv+2qejPAX0OrY2tB6vfIlRryV3mT4/bptyKAPds3o6jw77qHHgDUSob0EgqXj7Aln2Up/
E6/u8mPEmtzNjn74lvz8ohUbaVuRMQ1if2XgqRuWoKAYBHVz6anTdytS8lb9BoUUX0GC8VA2tdY/
PjEqGNfrT7gGvLqadjQb4+vIVBNeYFU1PN6cBkAWvIfBG80CXYuVIpl7jr6m9r8f8IqBIRs26oJg
s+5JkuY4Tm24XHkna3j+vdri57tXLFJY88qU6o+604LR81lUCXvqzqsi+dRJDQQW5lfgJf5hPNs6
jedyU7d+ojd83J70ZeYRxBtJL5QbwMMR+puhxPIxFqQNm/qH0RjPrPp1iWOIRcKE+v9OzMIHjA5O
3O40Q014RuJa1pSJSG3G+bEgq4XYOd4RvO8iLwsrwNBq1bN4bAcQJn4h6kE1qKow+0L94RF5usBp
DmU6xwYNtblM44e1U0VWoOlYM8K57Ik8Tc22OClTnwpnv51QCIoRKR++C74zzyVFNOTfhYEU8VNo
MhGqEg9XYX7prpdqGRdmy6Fzkx9vc1mgjxywO4msTN9NivxZm6xGtZ2z46X20bRWZRBZnP5OUpGZ
fswMFTV0yYI7wjdblp90chPLbol/gnDSr9E7rsluvQFYS2F4Qmt4k2O1uqGL4DQDCUG2cWDMVq+d
7Mlsc6GBf2IPTlQXrcJ5OKvgcfnxOqmShtZX1UJQ1OUOWdSkJ8WRTdwUb7hRRwL/zYbn76LfTGTh
F8/dP2bXB1UOJ6HKv7hzbSmkIaI+RJ2dRj8IeeNUCT3hDD7VKZx/vZK9RC1CEWlrQ6vMQTkwWhG4
yW4zJjYgInm/xE/ak//aPcRqRSoK4Vo/t8E6M70/2cZGlguj9s8fusQFnJzRHVEvCoFysuS4ic6x
K8ckiNT/W/Pm6eDyN4rYdV1Itv3Dh1ZCrtk6gb9GTku93ApPpLvKkyp0+YymLfkIjRb3sdxqibLp
qiyR/jT4On48hB5RcM91jwBdEvuq/AcvIFfJBtME1Sna80F8kqV9tkT1jEk+Kk6mREM1xJzxPQ5G
iC2SM/1HFl2/Pzfoln2eXXRus3rGArUFKUSLcxnqlR+Pcx+fPz6KOWAumfAv9oCqvQNPCgMQOcGs
r8U3Fk7XwGVGN1LzXWPVtvisPUWNtQVOj416a+OIz5SWEhqslbtNV4j0swwjWEHcAeRO/uD+qumZ
ZjmkE5bLJMFBo0rT1/zzj/y5R+BhfsuiIP6RAw/tUelz1qWjx7cDuiPP2ZvCSYHQ1ylSfniuFfCh
8dRJQhoFCdoyuNHptotglrt8/cOE8CqIDC11yl3NObOlnpGoOSBBZnz/7cqgLmkDVp3qikJDbTCD
eNiFN6OwXNqheCWj2ERmZRCWTq6n+mcyX27U+F9AHnNC9Yl0twxx2eJYs+uuCQTQ7YwoWbpmcVmU
iA17L2U6HxXWvXmUQAqmJdf9OIDLhe2D5+3kRftdAnpBrf9rM2muVAHPNf5qXhMaf4eNLpy0bojg
CCPTd5RhuZjGaRKMjRCY/kwpw1SF5dcfAAVqXG4e6FuVE1Q8FaV1Xy3BfaTw5i9gtB8KiBHipiud
OFURvzEEQxl+VDHkC5Y8zz0Xl0xj9tmECF9Oz3+qwA1aSbBaKm9GAke4oRS84PoLShQHrJLvwGEm
RbQPc2nfJaUMf34ROXwjgjncGQDuaOLjyNadGUoBHYeBhuqwMRgjrK0kmo63F67ZkQPmC6bfzHPQ
7giZi52tazxQezVKjkWddnWXuhEKktzEmfUpi1syehQatIjbCil/wsC0D7tU2Ygg2XXqA0CERQt1
JAzlB8GL3s2NEAA96OSMWst/sdt5hlqFLVgrPywQ6X85LNQAdOV5OX12qVL2mFeWOP64FvdoepYA
bBZPH9DnQFt+YshidRCInkcs1CEYNSunSIgYPjY6F2L7eNJ1RePlFRGABaA/LO+2bqys9iDybEDG
fjVcWf7KGlOdhLtScySGPawXoMfDfoSPdVM1ETdbb2cOPSbv/CwpvT/6AI00XqCo+LvnT61KBP+E
/i8lNJmM55Wy2cRdFSN6Gi+tL0amiSl3dt5jwbH+O5HKii+Xx7MWJwvTiECP99B2El0+sItlHRF5
gy0wRwoqrO1jqGYSu8unPb8qIA9LggxkpsMfRs4JfGJ9R5KZQLlWCNQE8Jcvm3xBmb2jP/JcioLD
nFYxQvsv53Fk5s4o6VtfOlAVdA0YlllszAT33uTEiZWxnzIx7VPhiib5wLRH7y+c3i/0TMgtxp6x
UN1SM/MovRY41UOMIpZjGAUaC3Lo0RGVLubWFxF57iUxaK/Svi3JxY28MYEn0cNT9RmNKSmbHujz
roy1KVH7YTxDCdcgG4Xi2TyrhlokLeR7MraOtLWYruL/oM/Oa9Vr0LcJ+UMU7c+297s1zIxYvpPR
d/mqLhhU2LMhMQe3iuzUNR60/hQJsJLEHGB8AYWiLme2LAdIglkYhR+LIVkA4VCOKsrIiSVhAATe
5MIVk4ONgDI8Km9LMS8bTaOsSw1SvgyV/d48m0pNzKCkB2f6pENr0WHXfkD/WphCra86qytTXM0g
M+TrtynrPqAXOxVVyN46b2bSdWi4cQGHUSjWEhRgp4D+ImRBnbS4kAiLe3c82TSHn7FXHaNX0KHG
wZe1YnXpsVdnrGnE8z2xVRogE6wCYMhcluQRxygHoSqD6XYOkDa6UIqaTec3gIw8WKkHXQwa+tGR
yVkT46jbR5Ou6+//tvfVsT4JyJkYlu0f7sBMTebD9vmtH5poJ836Y8C503gnYu43NSVmo/nPcD2z
da2hWRHHfDNqtYm5vWFPlpiOhdbgYHu1XQsujuC5HAEW0tpx1uD75Y5GnK61gJqW3Aj9wa6FMpEF
lkwfHFVBdMBzol8ZFpZVcmd6D5D34XhtcAnmYkmxoGIEoZ0v0B5Yt3R6UuaZofb2VAPTcLeC8jp5
shcYgqAqQOw0SEhkoudOQza2VtPd4VZlxPR58MOg1oRBzUbR1Y5iyHVdTlgE5RPdQCfTyfhnHbNN
7qcu7EBgrS8V/ViETXyw6kXPmZJyCSMAUwSMyczo82QpfLBB+sbskDY4agwKGI9ufSgGCC4FweKQ
EL1PCw21wkJpLFJEW9CjGDyFMX9mEFQlkFLlRTWf7XQkxfgekXdTB7Qsti0GtEvVkcVYk8/MVx4G
grw1qmeefRnTHEOFpDfjLOcjK8kGMD4VdoYxGslG7vljmP9osvk94JmC8nuYoHmUa7Ann4F0KHMO
yiK4lUJnjNHNHtm/fxGw4HFqSCRWPLjdGcXQ71qarSLMf2fwMW0Dj7fnDD3Vf4cvQFKg72zYnA7Y
utJw/EJdBvt5w9aE0A1kAoX8cRFAtA6wZ/vExWuVeisD+SOBpj3nUX6/H3LRlLsjy4q/PCliUNAB
SGuRTvJ3snjRF/6qaleX66qpKxNtdrDn6v1Vc+cdIW25Lk/SC6GQ/SImUA5ZPQ8h94aGO1pOD0UO
aBSKKToTLwMYsiCiAWsQYChxnkgh76kjJGffB4A87NnfBXn877Q/4tt+fj106izQn1nmSpIuR9Ml
WuTqr44h2lGIxTBi6bCRxFncdmQiZkMFFhxkSKs4I1SNpo7B5Hpk4XJ93bluQ+fuEjlvD/097ncT
KzHWNjRgwsyuJmWpEu9B+ej19JyFtNeJUdDj+/XAuajQG+hG2FPTJRTuFoL/4CaAtk66h1Rnyyi3
rURnEBD7b8ecPMS+il023flfOME0fD8eH3bFvElFu5pY86kFSefK2t0CGVcPtBzp5U8GGx+FedkS
wDT75Yzj4G46ej4J0Lu3z0mRogPdxItKjxqf6eXNNJDY4RPFbouE1IG5yRhRXGW0IByBxiRyrTLI
MpQ3NsoehB8Pb1cOxsiHIIEVJb+34BorNHw/LTmnKJ1IgNPG8+khV/1UfuUBYyFwZtRaSKtmLUq1
sYZejbar2Hb5Zuohe5ni+NT8OfSqb5yzhIZwvLwKoOElRwaDhHisUW3k/LuHRAbstbPErSPsMiXB
odjgvHz34/CfKBi8zN2aug+hBPkCdOaUxnZG1D7/Vg5DAOLAA4kIR0oeMdnVxQ5jtprSpnjvg/0P
TaanAEmhRCSvnBlM1WM+WHhtV1i/1HX7F7VucXdjb2A6HbvhGEfhR8Uz31qAy8KJivwt4HKWiuIe
UJcKsKM6JqDp24cgjSL9cAUfDjVBntfnua4ebk5ic5Wsb4gJcpQrrFNo/sOl2t9Yg7WYivmAnHnV
aNoVh6DKRuuTN1JhbzbEkz1rckJf3PHPjt5WLFCgWo5HCp0wOgW7UmROgZ32sjsFqaRXHBm9TRUA
3bMwhlQItu9oZfd/2YavIPGtMMiPCC84MVVCba3FaCwWfwBrKtBfmZuHp5a9l/tGbEhcrKoBOurl
A7BYnKmeLBFmPGHIpU4iztMuBiioE019iJV0HJ4mQJEw6kXeUOlXeDA4cjnQXTRl7cbaidV0rSMI
cbTG0zTu++K/0qusSKXi6fdpSnJINSoKB/L15RsWztWpaeGG/d0dTdKwL5Lacobie9IM2C3tG0FK
gOhfJjrHzy3tMwCSmm1o10mCM9PqorjR9TmFDb2yQjKiggdMsUY4wWMxPsyiUYzvylqHVBJxiP8O
DytY9f7R+SGcEhmbgVgNGVNqcZ2T/BNH/4fzaRuHH31nhHEt/8Q2L8FOTSvSL9hBaJIHaIixOqgB
wkYd6iCxZAJxTVJkTFbMZISmVEwycBRuXS5R3IV3fQTDDTfWbNBJYgAGrK7jASF+D3hylZfdMBbK
MuHz4+cVdeuyJ9EpBb1vcN0HV/tZCizwjpO+ILhAP8NzcLnIClDCNB26/9DmC+lT6nD7oF1+BPw5
PGUKfTCIBz6QfGjb1AL8asfm1V1oFa6JDlUdXthqIsg3Phuvbk0unrDr3kEA0Syah/h74Lx7d1fB
MfXqhMLj9mgaYXENiSf6xdt8RyshRjvUOYWNrKosBKg/eNeXXfhjTMGCM8WWwvFdy8ws1Mws3Kut
wrore9VfUfvyD/uhpLDYOLnAsxxoc7Ul7Uf+vsKCQwSpDc3gKjZYLS/pWDebcS8329BJ0Q7aUWZE
E6St40q7l6w7s+OmbnpI8ftlb6dDNMu8wJWBWQFIpaESXw3ijm5WM5u0HWvzUgDzW3YdmCIGEUmU
sH/AMd8nQ2MPqfpoqgC221a1mdWyD05OqN0AQPYKLKI6rHJeBk5FdDb8HNBwQiUc4xqA8kbbR7F5
2GbUt9L3uYrCtS+RPLXwU+hIOmyc/sXktrsGEDBetVXacdsPly1ZbqxLAPFJIDJZHYpYLDZImNDu
VzX9czNb+Z0FQ0eM5m+ZcL4oPc07I/DgTZc2I6TUoUBrlPNvDEMDRoKKiBxalirbHedMvI2msSCG
guanfKieRMV+hJpP7gXucNJbigfEXO3pAwKYBHWibU4DePPN2O+pUKMIG6w9JUeXzm1uLcrwTDdn
tWgBbSH3eD0QZixf50SS3NYZFAVnJ45A/4eFSWuHNdxRMCL53yLST0+4YIupe8VhxdgVTeyVP6h1
ypDTmZa5ovcP8U7Z+ORn7liRDEy8xP+sezF9aGLo7OZne1oaxhgl0X1YFbmBUbIuvW+djNiGDnWR
MsCgIqcnBtqc6jYjYejWyaOMKlQJGSEtAo4iTg4zRZ1WfPdEbccfCJxOtV5InjazRJ6ge19PRA4V
6pfcI49DKvsRByBVZ6B66DNDLeoTJRdrmt7ZkDQWINrGogTvUee5oYTx7rGHm66nPF/KC7qzfro0
0y72QCbKTh2F5YK0/1a3yGcg1yo1GyOhcTAr9SgMUoPtCD67sXVjboD3Bk6W4P/m9NTqSJIjaora
i1lsUCKtrF7WqCZRFis4DQBSs+IAOtsTza0DLUTkID/Jmx3mrsNoGXr+vcYUWc6ImB+UrjZx/XL5
guvrIZbpxMhcP4+AH5PZEalvEEUle+is1XfoJxAw7ydVLRVpsyCXoIlIcl03E3olctwXaMLsVyjb
hvH4USYauiGfJEYTyqgLIGfnWqncZ7u+lr63dQzVe/OzZHvbIOEnLD+nw627uvHDU2XjP+Ur0nIM
gnicKaLtSXIC39zPTEXbpI5RE3r72cGGtWpEBpR2ujioY77QmxSoP/6ErB6qnJVwiA3usJdZUTtr
UjlSSkzmsk52+lgTqqBVdAylslMFM/RYe3xoFfOtkBe/u6WB2SjeR0DEwVninj/Ew/ujzi+CkUc4
nuYIEo4yv2rE5zwMG9RvoQJ/SlJrlmEUaPqygRh+bDD5Yx/XmZiOSgzZUn0cg01W/VzOhFuzWqEt
hImzZJNbbmddGdRybeaURD9bDWFU9VDH5DNog3I2hZXgTYblMAdYPyjyEXpmZTyFaoFBqlu3wlpx
wxAMDOtdN0kP0bQ0hLYHmkpcWsCylEhR/uwyDeiIFg5W1gYVlgrwlH0J+8WozJDgsacJWWR/sq5d
0AmruOG/PJUQNeb6p02tGJlbHDXWQ8sF4guJ42/7OTJ5m9Fe38z6kopczouMtfdm7nf7h0lfTxGj
4lDobeyFIUeC88tzmLxIcouh5IU9fA9M+oMNVHQ0IzAKpd4APKAEcmK5cF7x/n4/XLHqIXn68gfm
Nb+1iclgT+eTcsSzefJbPrgIO7p3rAsnhVzrviBVnjRyTfKIvJ++GIoz9zmzP3haegHoYOzKaHCH
WhryntuxCN4kVkyros5ldGyFzEoCq/7AkgVj2+7J3JGjjfrP75pDDxHjLtWcjeAjuRHC+6CMRtrt
9rbXv1pOpOGmKj8+n3zZJuSdDkTMMu4qUiBGDN5s0Al5eNwWPyQONzY+gocyVcMFR0ebqjCBlukp
zNXM2/7u3nMiK8W5KMrRQ7WOUVXqOm2vmlYKmcTBB3Piqbo9tdDceoyYvx40BB/RWdfsBe3vojg1
Dtk8OpUjHR86tt7NCfJjlUtDmfRfN3ExJN5uybwpdfD8YIlHOQ3DQgCeZumWJ5IjQrtLX4PxFQPw
C35t57XdQIaHR7DREMEnwz2E6qAKiL7dBoB5e+aia/ukbCLKMD5pvQCDPHuPyOkAb8+8DOOqVFvQ
fjzm/8hBpCBT5F4rFaWOCUxKDWLc7a0R7M5rz4Sn5CfSJ5HDURutJiDH7TOgExe4cjJFLgPbIBY0
igEtHkpupQP0eQ7dORuhoe5nzvwBsqdpJ9EvUzfgDMRje0QmD782+Mow61pZ0wopl+qmbKEq978n
ec8vU65YbNE8Q55VlBYlKBgMN3StXU6wrYkSNL/IFMNB+bopEuYa8OaX81JDKEwvX5LcyL9HmRfT
ivGcBG3pgXnstD+gXoCLL6O3enQlJ0YVTs2gZoXAj9mbWMu06xBThp7Fyq2iKZlmPyMs17M5jf4z
42Jn12jb+C1SGkrCflfL9uaAi7xpdQIABXLiGnI4o2A7YQq3mr9q1BBq3ansdm0gSmum0XwHBDLJ
YKJXnt9vmAW5opgsv9HhSP9K5wSQyTfiVWPRAAPH1jJpT8jJTJ3N3WSP0ioCs83cokQvy28FDRRH
WdrkeE2t1wHV6o3YjgXkk73dr6BXe9pX5XwymXZ8zMVNNeJwp3EOpXu5FqFF0dm7NblgaXrim23s
fODtEAw7/rnStaLOORI0rluwOVvXcZE6H5J9JcDRPa78HeUfaBTxUcBWPJU6S1zrp9m3RKvdiWmz
ozAasBXI8ComLQclnGpUaSxPnrsvLn+O6P48VwonGZwO5l5PxP1K3LXlkXgz+PL2TrpNt8aXlJjZ
9qpMR18sVtsFMnjXEdeRXg/8Jlw3XctwNglkSJj19to+msk0HUFG5JYavMMvGlEqXd8fxa7Zobpr
CvcS8hfdSQYKfxWyN326pR5gd4lpQkytRznfVQf48I22WWZ/rq8gFf8MJ0H9XBsXSQu+8cX9a3uF
npHvOIEUbbT0jN+FMt3mBshAjYkrHwvlvW4nxUZDU2AzML5xlsremSKfg7kYd/bs7mIaf3MnwrCe
i6WTN7/Glhpb9Ye+RpOFuPP1sjhdi97AyAhIvDgZz3cxgljUGax+7oKdg95AyZlXKDPHOq9Rs5fY
aGDLvev8YWAl2OGgTnikQgrAVun+o6b+HcG0MlTz1auTmJs5abF8nuXqLTTugr79Tc+tZMZOAm1+
4XbuAACWMqY4MDtzSa5PkJlVxhM8fIMOh6A9sZywzb5YimCROeiWiIMJosfLMdqzl1eyQ3p3FIFp
3GL4SCl/kIJybGz6vpkOB64GCbWaAUtaWf1j3yOqyuuqduCYTvFBxmDN3wwHsGpd4CSYPW0TsC9E
HvhUjV+rg3EsaxgOH63/bcI+PDdMJS0ffHH6R3Ge5xm4aqsXmgzwix2GfuiOX2qbeTaoXQfH8D20
Tk4ucjGUs2BrXmGT1GP5PJzNaZUPh5sCFhwyprCvvKpf4ZOJ7vyt4J9dKFGDccTskvUyhgRmY9Bw
2lCDN9+/lahT4An/G3YQFuUNl/FtS3kbG3gy0HxbBOvhRIgqnABY2UpRxWrk7Dyxkp/Wt9x5/AAw
C0lUVEia9Sr62LKjjzOxk/uCgJ1S0DtSmEY1I8TB35xjRvAtvjmrA0jcjEFUAMSdxgnJVoBnB7ZA
3bPOFaCzD16uLThDMUrXoe3vuvERWk+Pj5kXgUuXHRkTYBWjexoCmzKxO6yipMEAn7OOis6gj2v8
KvnJXRh4uh/jMchBuZvTyV/VXKxO+yY7jBploi91td58CNTIH/m58rlFs0ifTKSrO68GI6lfOtiu
BK9HgNyaMyyjt+M6Te42KtSeZA5/fOAsjzuHbTdxQJtLmCRxywXg8gIHA+XK3Xmh14z4MAWZAAGa
cseS4RuF29BclHivwKezLtmhT+pPB1AeGdaXjSFTNurxuuay20mRqdkwTXZtjck/HhKm1eKGka5n
CBSJxikveMhxDBd64qLNnpQP8bR2TaslK87iEONuHsFc6HrHbUbb+55E8e/SvuwCaJBPbwGx5Tip
XuNPfB5bt8t8nHOj8wGNmTLjAnlrMtr0W0tUdzYLUadMA0kDKUSf+1FViQWrebPS6Zv2yDO1Xl+f
gDFdecjfK/TbLETPrs147XZvFd/i51UXAaVS7p7azdukaDEWTDnesYqxmgVgZQ2m9RADUx9o7xy4
n/bD3teldBgJmj36gZRBDKeOdY5auXA5V0HOSddzaizsrvNkTcFpn4U8SpRcY5iX3jEJkavRCBJO
UiHYb+HfhoWCxpdkKiMUQ2eEKdaCQ7Q1bbcDo+OS93TQvPCytvO3fU4yQ/UwmHc0y3+1Ylwafjrn
1xHyhHBhDChhEWMDdGYcn9W4EVmEhRc3svh5fJqyIXnSAibYWf2KmZDvtq/Y6cBXQMMapEAoFnrj
GtjGR1sl80sVSM+jB5t5xGnqONwTyV9R5jf0Z7hd8xVN+XhK1TmTigVMGIKCHJ+3urFaYcapaZ52
x/R2H9cQJFMhRdcA1jucIbGyPoacgDEhZX8RkHJCmv6KUE8jtEIPcjlx6kwU5AbavTaAA38Gxtgm
WAtALaIikHcPXFYRQQ6leb9kQ1lLdDfvDshT0v7hNKc2+UBIMRC2dF/gg1dFCNxx/zQfkTmgJCUa
YycKyuAHU4hp7BTC2Ji8df/eTY7A+bxss13MPHnlw2iyBenlBDXbwqeUPeHmVKkreH1OyJI1Tx+Z
tlTeV9lr/CTJ1MAn+bltOv3W8Q3qMDBJnGEuZyEQsQWlxCt6r3eXAFPU9qVDymZ45PXd1V6MjrPv
HbD+whJ00vzG2cbXR++aqoF062qmOupXc2/NYXJbPxHX2DBx5qt14ibmDcvYuzIXOwnQ0VGxiLoT
rQ0RxeivJvE1bSYM7bxF6XCT3URpLZ0h2Oue/5iVdDhR+/aMjE4UnXbrAar467h35AN2tmFGfmNF
Ep+1BuS2Jqhm+ypIR6SXFZW5w4IOYDVp3yLsfzAb3f7IlGSyfCrwBVWsZhoJcsGc0z4aDFXToW2J
7d8XNXyjLiHV+duY6nMA+u5h0oda/+hwIZpcNZTQPhbtNOnT7XXkjDZX5WLXMKVqbjxTZdfpfx2R
iDLGhCCRQxd7FfVw5l2p86x/QryfSQmu81810hi7HAKigB1v9yHAS55JbQFnA5QABbVltv/lJgwd
qk9zf4RTm+0ne8zraaJ6RVhgYrBCTDSkVMPoejw4m/aa9JTIbuc/t9LAcHsopZdUGPLxrXSUHHbW
TLlSc9JpfUSdDxCn65OXXsHBtKJZg2+GbJlAMFhysb6mCWdyl0l3klGO8aqqEpbwpk8IPUwbLSp2
0Sn8qI6eQ52Em0QJCwh8SJ2ZYs9fuyTTVPJrEKpjzXvLjm55QT/mHjOyuUtlYbpTBqPDhOZM0SZx
MFgrLhmiBm9Jd7dPaYdlJN5PsgBlEdB/JWtO01qmyfuYZoMb/FbD+oUSXcRGVBe4BNdPuNWzXcVm
uISiKFFATqcno2BEAS9vcH2adTUmQBJ50KID4CSVFdJg6IQYC3YxRir2opA1YugDgLNhImWBZMrF
SHeiHuBdDMnHEDZvqZz9tJYsmEAaDx9lIrzX869HV6S1et1pNXBRUcNEF6P89SES6MzRu4UTbju1
d3Zr9Wed18kEH8KMHuePA0Y5bU5Z8IDYjtpWFDE2vmPBGPix+o4tQ2mgjZ5YB79suZuRn3dTK1GM
EiOkVOc6b9I/E8SqOxxOWn2xXzt1JWXIp2dqGg7JEXJsroZ3CeuDI4q0dwp0iJYG6fUotioAz3ap
Yz7S6/MFFUBqcPL3CSc8R1naAHlScr70i+XZ5VaGLfpg19bmjqJkPyhI1HY3VICcRrgXWzs4by+/
U2GlwgYrJlo6eeDz+Pm8gN+RVurH0d6qbKPSGSFHIL6uyWj3+cHec8OfueMUY4nW1oAk9X6mSYtm
exq+8LB4RNDfzZBLVCcArp6VH6jipN+5z28bACxgM40lmlpTb9fUHEg0RKJHisYVI3rHuD9wV51p
GLlLJyXC4NLbWdlCFeBm0H+L1P+KRfBbk28Z5AE9/4PQJWqVMJ1X5LHFslIOzsU3aMFFR+inuLjJ
vhxxMk3RcRBVF4a6Biarc78Z3KC3NgbEmaB+xAThemdzpNR/Yybw6kB8alg6jqY3lxxu7phuNrOK
E9J9c1XHVexgfaUyppr0wVMAt2C+ShKDyh16uUU/sva5zgUHJ1D7q75A+WyxO2rGNX01oE68UQJS
LfUhb6xNTmuvR5z8K3k4ZTrtWnr/TaZ6OJKHEW3VVpb9iVaj8xZEqpmtwsLMCNUmRFVxy6b2JiF/
S/zI+t2g5VeVR2X7hsbLj3capms4umc1nL1EdSHm+c7Ju75YVglbIsjhVY6y8ZhoP4d3ljooL0OE
CqLOs1m/Ixk/EQDbsQzKW9KmTJC2Vq3REXFHOH1fiV7eQvHb6ShXf55mSEcTeTgKzueRld7iK4O5
xUzMXPhEkBmwf7jdNeFE34JwbzotnEK0zP82lWxcTam3U7t/pI6r4R377VXqaVA8le/YPHYwOnJX
UPV5jjSKDXGwwAUeHLc3rvDOBF169/d9WBiswzR9H3VlbewTZLvqbZ/ki59jxzMEdU+cVXqVBtWw
VSEaL4NZG916N8MQCSvGnpEewYvnfc2SLeWey030/TcZDxI8FVhjU1cjsy0TZoH1wUWOf25W+ifb
hwop6dtTWFt5Mv69iLwPk/ESnLrBOrRNFfnhine+92UoFV6FyT0tZiWKXpS6flpiUP1dlvIb2rQk
WKnRnD/dXkhpJe/JS5Bedl2AOp4Mml1HL5SMdTC78xn06yP0vUqI6nPWUAJCIIjicRLfeUljy1p1
2KRv/zOzasx3rQKbaJvcBhs4qB048kjybqgTfHKVjEdSOkYF0RsrlwI97Udt/+jLZrqHSRLcHEKf
VR0A+uWFLHyhRK/p5F+ta/DwZYVeZnPKek4qSxRTb7fa4/vscTwOJ137gYatJjKDQnyJ/gE+OEci
L7SDWi6DArDoIlTAF+gzOjoVH28hKlB48w5HNqaJt1G473P/8y9CT6fI9c4BTkpzGx5bO8Z5E+U4
VAhoNVmNraPY8yQJiT3Ts0oCzf/RaRZbOhJqZIkiW8cqc5EzG4c/SsLfCMx0k8ENzBWLYkQ2Ff37
CRULIm8nfoWPdpCukgyzdQENGaEFAYHCMm697naZnlmwRBoOXOiCKoHSNz/9OcPf8XKsxLwo3H0E
0w6p4/HRG9fWWcce4Y/8V08UxEY+THwZGaGagnebj0WywicmqduJRG6V/zwvHlX9n0d+t08RuXJf
8vjgZSmCcDLRiHUdWJc1J1z07MZE55xxXDBG2PjA15HC2Eh3RE7PbPJQNSbkNyOpffwwmEcQn/6T
FlYu+GSYGOPmn1wNW6H3lcEkdVlpNYyIaQxHxe5fUZxhZiIWI+V3TBtVGN2I+sH3zL9l3SqvYZGS
72xtEfFcVPsJVKUSr3O/sIGHhCHYqfxi49EmbcY3NfSi2vZFc3g/gyUVYLdp1V5lmPUlyEVR6CBi
7arArxbDmLxx35nQNOxNn6m9FEFMNlYTZj4BxVJ22QpkvWiJGMaXYqJm0VS+7IHsfo7HJ7WRQiUj
++sqd9kqr8t7DKeK90WF93Grxs9Fwi6kIewDDCi+tvm1NbC6LThbYbEGY7+jK7r2SdQQLFOaI8kn
mT15MLy7sSeM7+xBdyWgtXRkoSMC43KLM+OQNO461ObvGZbHIEEVOv8MMAT43X2li0+iR+Ocj3rE
aR3B+dbOzEQoCZgp1+6S3AUyoTkMPX4DuXmKdyATVioBNoAZJB5mItvxg1H30zaizsJuKPZp+yKA
icb0faXhVm5iHv8Aw/fgZWCIeA7h6ySJKYmYMR5w1+A1orjEpqMWdqETVGQqdpd2kVYqSnlrTvuB
Md4RBdJRQAUidbr/JfQ7CAkF1z21NgnwApeW9FRZKvGbns22UsGZlcgK9O8hzUGkD7tK8iEnkUtb
eHd48P+wNseHJbN5dpUk77Ulea+LYsHbq3B2ceCY4ulpHCYEc/azyxB7zSa0obmx3D+uNZXZRPUE
TiwZXggs/glyPB/QpmngwTgSf4qTxRnyA9nZl7gf4ESRRWh5k5ReOb+UCEBrRik1NMeWbf+r+q0L
4rX+Pt6NBmTYtUtmFDU+Iz1GlHSPYJ8QNOqrUqy3U2rvJFAlKHZvh4/JL/SMl+cRoKieoewuHn0K
GsNYUeXZvdGMseO2gx+V/6zLJ3x6Dgpao+DTQJ8flwOsY+q+oClsOOHgl/L48jRMQOIw3OyNZks4
zg5kaGQAOIJYWpjHOv/Rp2kt0s6RGr+LTLpbXePRH50AyBGT/KY0pzrC7ML9gjzolkCBaKROS/lw
w3SmJDVplfKKFLlcg7AiGVhHrHOzxC0qw4wcm3qz3CCSLoCulJak5iFTn51cUuzPk6B8CUKjw1tL
vlAnj2DT8MNlJO+Bkhm+mqlYP8kwm3z+OzKS7LsCsCHjVmeJ8Ut/XHuxkOizK8QB+ldvLcrbCwhe
Ojl6QNdwNoMdCJ0WZXJ2+9r4P9RHYPe9I0aKYv0QMZe05Np1E3+KBoJgsyi6J+kW0/yBZvk9+9Q0
13QoUcgRF2QaZT7UmHXINpdY4JWLGmYgZtHtvJiy9QjOoIxX7WVydckZAWIUEBKmpj55n7B+EBJ2
RDNuk9tl31otqtZlOCXXFGrGT8h034aVyUNS5JA4DeKqjRky+HWcLEqh/RzvsRcc5FpmtlRkNHCR
xudbZn7n81R7UhmvmxgmTY64eSyXUCPuhMOWqoIMfDAeU/M+oMe1Ihd+DehSr0egdwkNFbn2vei0
IgW4/bcbr9L1jZaACMARhh9KAhD/SYfsGeVHrSbOOFvHrfDDOQM79aO+xtnNV9qd9anmH2ANIzhx
ZkzMvlCGUZh/4MbNWFctWPTODmWCLdtKah3oaJeBQFtWjrjSg3Ph6eKPyZ/rWOm11kWS3WSVswRz
Al9L6jI4vpU2bCH8LA0AXMS0AAFUPcuk2vpgYAzLDhxtIKCi9zxvjZVVAaXaw/6EIlQhcQDA8SCn
CpaKLwKdlb898tG+yqj51ayXuluIp75lGHbvC5JLdkhH2+6ElCIEJdTtNfnuankPQlCDMsGIVGL7
xQguDXDrSOJFnzyxBfHFZqSkyMOtbuIP6cBgsurhT4mDSSMVMWWLy7RWjnHq2jSiRMwmcc+V4+cY
ZMAbGeDeDmviK87jW3X4lCliMB54fsoAQKdoFp/igsTdCnSm0EkM79Yuvtao7lkzDB1NdSUq5rMO
0p0wtY7klc4gHBiK/8IMHdtFHyPM/OVlAMG9mc9zYC+hWW4b3y4bKQ5myrrMfdLqjbMA+wbUqL3K
gzwhoZn8ppbVs/Ipcxa7JLmcX6H6SlLM/UoAujFBAVkNVy/nMUH/JSeoHnKZlRIfq/T4iSHHc/Zv
+UiPXcsYawdIMdy4ngfNqt061RQGxPGRTQXcbohsXfTSt3ep+0Pdf2RpvnarGLBa+OmbVLt8R76y
kv+2MXB8f8FdlCntJDHxuSvGvG3JwGaw7fTDiwaPDAxY1jYEgsPKwO2XkNr2mK9vBMHwgOIOw5Kq
fw3MV9mgKykFVnXQmDfgT9lsEV4dwdPoW14oBmq72LkSi4Er8L+PEwsNOOB7tO7T3Wu2XgUvNlra
aCDYw7c+Tjx/ErkMaOP4GPpISIu0mC8tsw4uSqC//FNVDouMzna6o0qbknjogVARaR+LUvGi/DFt
xloLmmyqzuDPpdu+tT/O7DpF/u6vLemkekoqRlzSNu2NtdKqnS3Qzvsrr7WfasVpPQ1HhhadCj46
7vKtogfnLe2bcSmJfZ5tpnXMYfcKfDiiuNk26oshI3nYh0/UOSp3c+ULgDIocYLYoQCud7DIrA+L
XVardO59xKAqFZF/6e2OGE2vZf6f1C66zv01QwhC1mPSWxTtEcdVCQYNkQw+UOpHRHnNm6CDJEnl
ETL3J6LwS5qKutglQhVtTIetxo/VyO3LtD9wx2wCzlHCq7yEnq2HA7ReDmFPQZUyC9K3fABGJjGo
C591hWkqvYMjXXkavtgf70w+rH+2C7AIg4MoUEr/v8+AEnOEF582lFwEZMcSA/5o51rDRGS/DvgO
HouXWA/F9Q2hobwkJrdh/qGYA7qBAN2Qr0KR5talmQMReCkXxfjyOAxL/8Rj5xkLv37IBdsaMpZa
CA015OUDgAc4jKuds0SE19d+IfWk6EV+dd9kMN1jJEBbPpHBlEIU9/Rl9sRWlCU+qRbvDiB0UDCI
y2W3/pokaFQU6ajKqP4nyegvtGiHQucJs9v2uq6jmDpdLnNdGgMnGAS1sewpuKaxx7XVfjOWEDsH
3jLerIgqbUS67isKK+T238cZQ5ilt19GR2MtD4LNL3QLXVUsFw8ZDF8igPlT1GlLh4PE1KgB308E
4pEQhvmREBpLCeW//pUf1NcE2vOiKWZ3pNN1yCtmOGh62iL3txy37653mPbMnQssM58jXaxFlHRO
1ePiWYugxmmfEunrUTBk6WegryULCbLujuolpYZdL2Cvr919ao6jtK9doklAsu78OWT7Sm39M9aC
MtyMW+jff5WLAjbwndTt1rwq7jJiZB26MtJNHKq3yl6zYfg8HC8KYwI+oJNQDepBkelyg7bdjr/R
EpdhVlFj4hfCR8DSIscMb8Xnc2jZ1h+X5rR4Kqm7yfET5e5dsFHtxXBYC+Vni981338Wn3XjXROL
GMIyaJLbOQfGflJDoOkn3Y4vJyAczw6cG/fE+b+MrMsnUxsFtsZf2L0gsh6ke/gFQfHt1JbRIWIx
K7WvLutBXBo+HVSF9YLQBgpjqfumjTLYiSeX7DsFko6QXgaOasHsYkmto3d63XJM3n3+p1ikAG7Q
5kW781tFoqUssyGC1MR1O763Pw6BcU1Zz9bBY81654O5zOKMoQbuttn4dspzQYla3QD5rGblzM5P
ABkwpeW29e2S3bihCisKQG3S/1BZgQpfpwTRvojTK4RA0ndlfkVx/2CKIN00q65EZXTVKSWrjUOt
bluqfcyUzWFm/5qf8YW3/5xGYnIXw0cG2dOM8rwX1HVq2j9z0ACTQr4HzZwdIH3v78joLBl/W0LQ
dGR18/QHqmRI41d2I7TyTw5dupNegZUidjJzyL/vY29CggRHuGHHn4nXrg5CUxE7OeoeaN4zIf9y
qTPP3NyNR9vcInXEEIPwezCtzbRPa3RZrGCdAVt9ng0mNrXKyp+eBiV+s1Irqlj7nM9tet56zzYP
txN4aVM7yXMGBfhMuI7mrbSBvYhfhmx9RC1y7OZbIlOu+09dchOEjXan/jAQRA9DgdY/hQ3RcjxL
97nWhosEm11QmWV7MjIDntKBm2GFmMkvopvGzgamwS5MbN129zfenQMDkIGkWvBD2oA/tZ5JklPV
wIuAyuRXiCTZKCi+idfee+WOOuT7gvTfHUNFyFRpxV+M6d8f5qPDq7SAjdN7gC7ud69L5CnpfoYV
BIsz8fzlwwI/9oJw7EurPdYpiEpo6NEtaW4nhiNDSaSxPnJeri2kwzKiAkg/5Hlbxf5F6bmYnXrA
TvMNY84gngVvPvRWp0FkQ2GFo90qvZAGX0Kbm07nGtcE5FeikNGnazO158JnsNYbqYgqBoPpNeBv
qf32MdCpeqmQGjxH3Q1SYbgRRMSpDcIVWzcmR56fIApXRI6dk5WBBbYmQNGbpdSg1CfMMMc44e4D
gl9PFhIxY2MBonTr2qhPJkle6jfbBGDU1caSEPaaMZnMZEzpm0XzSonDLAvsPk1/XWdsSebBVRII
x/97JdbawWb/9zhwio1nnW2NBx+jjZ6PKuu90oumadqGhOiZd/46/JTcrdE2Lmx4f+I23m9vNFRj
bzErqPgtSsBDNznvfOIbEe22BvUm7A3MXKaIXnn1qCNTESkwkqxMl4L2H3S2YJ20ZoHkGNU0zGL4
D7l8GRi+9wmUGZVR7VpoU1oyFodn68D60VnIBVxig3LLogK0Ir3BNvOZGwmviTDW6EAYKbJkE1hE
5XGf4Xo6o7gdzHmB6epOmhmc5sYrM9Utis8GUrWqneO544wMz7Lnzi1zKmaftZEqU5EMkxzPvGhE
R2xR8hIYJ1BKVSdRfLks1BCCvhezNQk5dXBCf7db781mOrx2uQRp5YHwlPjiD3xkCBUK72CIKGn2
3P+dwQOxQqsJbxb0VS0otiGW14/PvxLzyJ1A9xJbyjsoPpGANJXdxe+2oOM/akaZ7vMYdZ08/yPS
e2tpKu/kPQoTUneqoMVPTh9gNaHe2OZCv3N1EX/VeGF9AOt9PEps3eNF5plEP0GKI8M3sENL3sfL
79Ua8x+L00jtEqoA91ynZWTZ16NLzzoxEKmWZtJA9QChlfAaPkYfGBIWvqr+SLtdflmYBF7qfQfj
BaeMYYVFvPd8j1w4pB30YzuryMYXijBtABInhfxJLcVEV69AeSYv+Ojhi+ypuXjPhClC9SaZCZYF
EdGLqaUZXZeBsPsF0NNSms9PuiNzx0kr/wp9TcifasnG4GxkC8arOTxiGng0nXYJJrKi42DO/isn
txg2k0oZfvBwfOl+Cuwk+jRN2FzYRHRgEYOW1rjLozk0pRYbNV1rublLusZGpi1R0fnpfx8kmlRq
viYma7APINoBPaH91fb4mi7kFFC8gKA8e0PBp2CkEF+FyzmmGbfDqIxjlVN7naQHeFCopwaeNtC8
rDjZGIsp9KcPmG5wEJxl0bDH39+OlGSa1uvCPPk3wRgDG//Cj0eCktniQ35lfGTmVZ04Eb2bB6cK
o8lHkrnwFouP4EqFCJXKMN0aAC4VWcZq9HG8FaX71vBgErlQcDsTU4pzbKIePgAmaw/VV0ppRHBi
aTdpDg0QqaOlUQBgEW1oHd+Un/jAmm2npMZGuJXJ+9racGcTtmRG7Na812zRod6XLwe7+cVD4hhD
rQcmXQnDxkl4YOgpl5Jes16fBKugSNRJPHLnBvId5alNUBG40TmWmLxPMUeRKOKx7WFVCUodTIhb
DxRo8dPbhm0r0z6R5fUpN3iWlp9o+pBsFDqMcbBvMKrxug9rriwokA0UoRSwAxgrwAvyU4t3AwFs
sDPWWC5XtlAW7OHzQmuRBb4nEFp3XDujFAHzT0nqACsB1qJZVlt3nnOa2NSA/krB1poLisgXd+0v
1NKWE2B/ARquv3RFVYxoEtdZBT1ZdsKRCam2LFjxX3e+p7J8jQ79UljUMjUswiFQWejYHe70dISU
i9GszfVLJj1KD72Hsq+OGX+WdyYWp/z5F8joqFaHBqMmgflUMhSmXwod6B0IO/dXkUF7XB0txnJz
KY6o/JR3UTB1V2e42D9903dteAAhCQCljEX0Zbd6l9uDYy7RS9Klxy8T55UAph8Sw6b5YsnNyKwl
QHUEjBV/n8u1mxvL14l1/c2qSDv9/UlPQsPAp/T/G4Mu85nes6NVg7M2FFFQli1IzIski5hhokr8
2i642MqSx+EmOA8NSgKd4Aeg/qcTC+4Dcm9LSbamdYUOn0+VWd9yH87IDr+A+BUllPo9ai4KB84n
F+3nzL58AuS0sqYRXwCm5RcjpPMemNZNaK9qwLJkxbZCEoQrIfPqfyxQ+v6f6ZP1yh56Dcdh9S84
nMA/t6FsLCgRJTUx8dHWvAX+XlJq7A210BGPdlDULijnxPm59pphfCanbsq5kISUkW9azbeIV7Y1
0RENuwT7E6keDvSe9IwRXSjiwiz5eqtB3Z+8jY7ZEcMpdZovULs/lXClaxxGxnkm1910ryIGS0hW
6Bn1O4vJWfpTNEm7UtjlCoQY7U1RxZPIQxnjLLC4k1pnL+0EEnAALSJo+ByiIvQS6+poEVpdR02Z
AU/6UgDaTwbSFLrqFWaSyUO4/nUFYmsBhrXRnY5T3Dc6JWRYQxj4VM6GZohh4ybiyUazx6pwMsKV
hSn1B1kPXiw7fhkhMLIuq7lAjNbavWoz9z15gHq6/RiZb4fx9EkxBHfvfCmxi8HHxOgR2k20aKVA
PMeDYCF+XU4yPjMo5Zx/ukRVW9Ya9VMql7HWudDJUHAtw27oYXEZeAX6nCwsYLvXcCsKS6BqyIvf
YevOsQX1ZNGvX5lDBHmMwIKf7fcLjNDb+vXDuEYMo0TIYYf/K9jCxKzJ/PTHMCEApx7Tfr1K+zvu
bcByAAGrdfzakvjyUNpVKH9tCiyuxezMnWlxe1t0crEZlfXPCElVJYoy0hjdbqWgXiFvBlBsKY6x
NdnUyp04JM1TE1gvsdPqKIgX8hgvOmUsihC4D4smyzue8VTNSbOyZ1nUUJK1vX/4pDldOSr/YRAQ
sT6EtlvRveCkoWWahFHx75BQhzm/tXvGzhrqQ0kZJjZWLi2E968ohm4T6wJQPb4sm8T2b/1WetAV
YXXpqIbAcJ+o5rVL3yX66TpPNJOyeeiB4AcSdqhjQ7o/lpQ6mBpTzPUu07WYOt2xefye6fYjk9uz
ydSSKPlz4PDKVRK+o2QvhuguDphXZ5Fk6dDT+wbRafQLZRKcxz2CMbixeuculgzq1ok5UlXbT7lN
xJDa7bMlrfQ95hbYBn6J71AIB0XIZKS6rv6tUu5smwPSh0T8IzCOsso5FId3w0mU+pT6miLHQHAz
BIHKTeyrK9UEpZ2dDXAgSLxDrWjRM0fFzyqahH0STIMIgiTJmXeHdNjwpdUjLQUwgi9CqvQSKXMP
HKoGbwFCCkrr0ehef7fahmBh8IDIj1kaKavczXaCszd7zDvHet6E1g+zCVt6yS4eGdzzI2UV6b4j
6qMNEry4rBCMHVHSRangHLk0YI+lxE2h27yhLF5bdnXsGKC8FfU8vOAMBf6zd7ufQC8iig7iwf0j
/t1lho1IfjfX/0OHBH9hsb+1bD/Wyb9whONeagpUDv8GJ74sQSZ1G8HKjeawXz7ayZwXfsyWBDf8
ZC9cPlhAI8h4dnOLBAsLdSFywEdDkuX3Wca9Zq2rxq8gL6n4GUxIBzmjmzb+ckQbZoxIIFYhkqcK
1/Hz8ke9/3ZCrKSlYQshLs9YV1gFluJA34kDW0qqUbGg+a2aOcWJOukNQ7idX8izL4LSn0951qST
PRNV4HE7PhKEMr7lZiO0UwB8FxsQPl5J/x9C5JG0BILnv+NapN/x5iveh9Pxoc+6gUSATTf3wDVZ
5Pq090MQEKPTXZsaL/IlckZ1eUETcWDrTc4VaGrvNqr+a1S1jzHLukLeWHJTC20C8sDrujvlGDxq
7CrrDN1hONDcXHaTgV9xmN9Yy4QfmsPATsbpYrrUiTMnMLAZCwNnJ/jekTI6Lzgd2i2kfTrjue4/
OV8wDnPdFC6qiikQChwipTZnM6JACrFjljByWy80o8SZ1JRJLExKAZHtxTaMb1r7/ZM6phw9CkK3
WwHJUFmlvEFlZyqmQwr14iR9zHlbhLOLYvmW+13/s+cG2Gq+c9ubLimdv7w5u9tPizIOKU8dR0r8
BEfWlSWMZQBo0XfmAEJuO8CKyYvjicyzqMNz8noBCBq0M+psZ9UjkG0BaMeiGdNYz0X3CIs7/2Wd
79Mm4YLu4lPS5oLAv2HyCRX+oDYGCICDfJq92DZmu8so/rWcujrtLHjyenXK6ThIP8+STFaNLZsw
dcm3HuBnnDE3bYhE5c7LsyeE6duPZPfi5xBUGIIhjun/O/kyVu3Ajg2er68PyvciJzCtfbjfjudl
mIClSvGAvHJn5OcHUVGQ+q4tBUeJL3Lp000R6RnpZX0mOIBS1ENTrvbwTLAjBOIsUG4FpB/AV3ED
+36gZCWdIuXZoaHKrls80ND7ilgyXE8j1hFVVsH82SvE+/FFoOFJZnfoYKmmGDTgyu/x/wpn9J5K
uUNlhRf+mrxdbtFOSV49YPHFZCxm0acnZuoVNSourxDUce5xjuOY7zOFGC0sMrw5mmN+mtw9dJ9L
Y1MTuoTIeVEAjM0LUqpwccVhTixeqdnGMdS7+AGAR7gSZfquUqOf7/+zZPBbWb3LRYI2Jt31Ytdg
fZbija2ma8W1POWDHMdz6qXDVSV0nFDC85HVxdUgLSh64KV6BY6Yv5V/lC7lAWwpK8JQdhmEAzLz
aeZDbsufZtAG5nNjQaDkxL+ccXvZx6Cy2hTn+f95veHFzL8dYRRbQlm56Yrwfe7dYZzKi+mF6rGi
3ddcrC/yhq8ny4853SdDCNIXkOKGw52zrAD3PilaE9Zu1g6ErhcTYD9l192lqQjNiZQcJ8Byp55b
tsfolCWgZ3W0A0G6c8RQAFO+ZPOXlcNdsUeENj49DKBt5j5uFSeWzfyFsCOqWchInbeQdhYl+fpa
nzg4u2Fw/Oz+RWVbcutARYT3wQhYuVn67ABGXqFyptd9GWsVK52ubQSISRa42PVfe+07Pbcv3F79
ZAZBV1R5RKKm2eroZ9TuuatIKIP9YLkKYjp3DTpvWPHdIncV1+8vz4W8zbLA20OxQKoY8JxLp9Io
UyIHURIJn5yP2NoWNjQjx+sjjvtxsR9dDLEGd5/7xXhSMiAEl07iz5d5ES5W/4h5Y7znws8SPodR
TVAay2CihszxuFWfFsiR2NTfXYnpO0kSOH862K2uR8NrGUgdTOyoXjWl+a4Yhiwz3ssRcLT0Wqri
yWzCZvYKEX3Fqw2ZeU1NGwhSuKOTC97ytgvD/WkWO/Ol6e+JmDAEZRps96Vs/T0ECfVnxZy+vfqg
8KFGlgjn3Mn531esXJTTs5r4o/p3ABfH2b7/nMZCInyULKMBZJbf/nkzQwQM/FTLfLy2ETQX5S/S
S8zGWvGK4MovSnQwYntjnrNBdKsKTXiq3rgG/ZPSd7+9jgSIdSwPsyZ+UWTw1Q30MHK3KPjAWC5i
aBm9sUcraSSJPq0KWoWMmYZMNq5HE9nqQtouCOqPJUPClsLZyg1kTOe/RDhapAIi7LczdUvJwFUs
dK8JHHYTZImwmRG+xQ/tmeXdJUNoh8oJEtO0bfpVTayba84HatqhLMhkjnI0b1cAUcDPW2SPv7ue
BFDzedtfnZsqzshu13bQ4F6nEMUitHBqGJXfPPgw7EpYxKAgm/XIECpWZkoC6/wurW/schNG7Uio
vMmXhecORz5jPZu+5STHkelUvlmbx8iLIH95lbYSYfGvTyum1WrFGNjoeW40FGJn9jFcBSZv0uvX
nP//vz/M98VPDbln7dmuIrH5HZ6hFBej8GuvF7bu0UXjU6W48Z6ioDfQCDMsdUfkf17DXpugT6nY
0SLKgHLNh071i54qCw+1/sQWGFzeN4qCvhbbwVlCY2cvr0mf4QeL62ebTnyQuhYjqpE974lOT+uo
St8cLMA+b7+2i/OcEOp2oeAoscER11zvUFwr6Y8RLpxklej2qj4MRcqUEL7e+BKUzgmCSIy0+sLP
M9qEn4zgX4hNFk235h42qgxY+in5SLLLEcopbfR3oZU//4ODnOaCwxRUuFCreFoafgsMtNHyNOS5
8CUz0OFv+ar1eofF7rVz/cpFWw0OJYmlRaE35V1+vqPsTZQsv3lkfhms5Vx/jkYrxmeuXDL2DV39
TVArKXrqXcCTsLpH6oO3ChyA14rpy9hEHbYHur3ucASsldzhbzZUFXptcEMR0Oab1a+8iF0MpTfY
IaFGeFlDHyrSRy+DsfKFlWl3S6IM6BC1TS0ZmWNuu5Fl459Rzxm+aGvfAVdzs4UXr2D6IrpOgk29
zcf2LAcyyf2Bl+ZykcZmcx9OOrBT4tygRbLofBodxwzAxVflNwMcWh1xaE7qmuG0GQHUDG7dEmG6
Kc+5VmAe+hfh4T8VBXLXB9iNCBiJp7B0Pt3afAY1mGG+YCg27Jk01P0ehIIKUgpK69uWRQY1mcy3
kGR1JAQKfz32PwDQQYYk7vVPe8KJvf5+Vp7ORf+WjA0zxTWpek5oJSDC6j8XFpuANhd77TIK2hSK
RS6a3+LNQD5N7n4rZIC/muPOqwyMQDoEAaNIsBCa5owjW9/j6Zev4aiUjwfIZb8f+KcUwHwBIJg2
5PS515LBLb9piSNnWXla+ARndHQABjByP7Kn8w55zV4NZiXkwDt7Ddsn/5ZMzZs6Fk/xuyHzv42v
Qmcj8XA4Hcqyxek0o8/mVOjQrvlwnuEjwPew9+vdNHYJC/Uz/D8XfUW9qaNG97c3aHyZejJcgCgE
ROHlekBSJAML8rvQ1ebvtLc/v013116ebWIJXqSeGC0JDIr+0WE5AlLbE/cxMTWJJSAI24eZ0pnt
xyCrpl6A7GueCAttzsYIjPH0MLLuCBfm+vWgpsT+DupX7XZ0HW1EHyOmSC1FIWr+WxKudLt0Lwa/
m7V1xXiAtk0fHgk9V53Aq2560JdIWJAJ4OzS1TPGWQ2LuFyu04Rh6d9qpGMsoJ8PWUp4YqUocR/1
+X4F3veE39iewMiufYFzVXUGFWLc74JaSXpVDpTbwpasj/KbmgH3Cr5TZzRmPnLRb9J/Uw8X7azl
5xgr4HdlC2vgOnpXS1nlhAgnmW6lMyPWEoHXkTaeN4sk1NL92MeFd66kDUv8DTqWbVVHs/bYdI/x
nLqLF+JNjjejsmL6cL2mRKZN/3bgRTyuCSQupOfGe1eR8gF2KIrTPojlPZmkJOJFKyFN+5tM/7vZ
4SU98fDsmfaEB6TcE9xgFHOee7hJ2ztkUfB9W+2/lXBqyCDGY7IdmzVCO8b+lngrgwmKT8OVa0OQ
PIGxj692tu3FR/NxftK2fBmBVZO4rTPS55IDEAoEmTRNQvJh9CC53Ys/12nlYBYHzhAW0mjbuuLW
0zLt7k9NiwTCmKen2Vt5zScQTJAUUbjoO3HFeUp9WuqHPwnLkWw4ggF3EN7XEVeizJpo6Vv+OiAt
50GC03xhj270hp5g8EwADL7i9Sb5BeBoCXL8TRzTiZbH1bKfgIbaJ29/1j/6ZyVaZ3M1OVrAa2TL
P3/VlYgH3kryeldCSk+3WRfgRPVsuBesPcuWZWpzveg5+inpQ+ZJO4QVTZd9G8G3RTJ+VMg3kYjN
LNQVnnuD4coNwakDf8h+ACWLMJVoe28mRfEC3DGKT64IIkaHo2mcTdhFURPSFOQ2ylCXIsbDeCU6
gzc0OqvcNvQ8FpPguHR/Yzhw0ppUdsaHA03maeomhBSomD3j1AZZ3aZiFUjpjtqak96uFI0OXwur
JOBjEUYVcJ9JiVLK5wxtV2vxxWgMuS9T2QHG5UDPXTE8vQscMmSd2VdWY16bSWAydylzGi/8N5c7
VYhXjf4NANrFVFidwja8KBpqGBJrAMVuIJO0QioRxo4J67eUjyXZ2p2AHXPFDYgmlok3g7EwQf45
EXaZAlQ7YB/NZKyH431/J2FCU0owp53qjaqPlWvJDSx/z+qoGzzmwAkeb+inea1+ig5bMAeNDCSC
4maV6WVtugnnE5TNt48kCRb32VCnP9eZhWT9IU3UzwI8cFTufRWyd2D0jdYybELDM+aDX1b7FtKj
JKQyEjhMnsAtTGYzJxec9oUGx0Zone5J2oWeYmnPgl8t+LihIMsXMQRdsVM8tAIZXUmwrSXKHMN7
xcW5HOmAeciMAIqVkv8ZqaF15SE5pNM2YM9iFixb2SDfDFpt7uMcumuLj57z6Pq1Y9si3/jJQ4vY
c+SMrvfMHDy3nnadZLohgjJBrjT4MqQlFiE+YioRclBOBq/aeq3QA+qBZlMY1d0vMB0h7L3Ahvd2
zWi40dKz9L+EbQuAErlfIRCCtw+UR1jICL1bLRUaAB5TaKLAZIER10KqlNsLA7qrZre9rpoZxmZV
GRQWdcbbwKR2TEtJ96gSe+ENXo4xibPDt34X3+5O8KYz/E/GWT5j9Hk2Rpk2TOjEiG+0wAK58svn
EsT9Pv/b5QRj6G04ZzswAdTaRmEt/uM0OdTl+IQFiXSYSX8GTayYL4KnDezjLlFqLfZK5hf2m4Ic
BMM8Mi6tImtq7zB9H/YGhkeqnsCXlLElNMomGYMSD0QGBqD9Gf98SolVh1JhSxwtuXurcu5ir0k9
skuxrirQV5dr1a51fg9tqSritarLvcsStnFFHiFRg3m7GsAXzecUhiubr06XgK9Mw2j/+sgmxqYQ
9XCSgl/KvIISFJE+3b94YSTbss40eta8x3ZuJSwRxoWdcuirx7S99QQ5ZTNxMIl0W5ykuSNMH/x0
9QoX25opcwXQP9Pn74Etcc5NcI4wo6s4FLxSbxpN0E/ebq2wJAzc1D1FwLE/6nRtj5mt8+XKjB8E
8rd0aT65C6Z/ae0B6287maur1PuoSRkSH9QkH7z3cjt1gnlP5bzrEZY9ac+BM6Z14Zzr7GQ6wuTm
C2N/8G27Vo/iiQH0G7I2l5N9NI8bzw/epWOvLDGytyntOTroNxDW8iSrXwW/Sb2JcQ8D9WhVtffD
gVrdqwz2mIyQnM1QQDb9yxAJn8xyK/JNcducgugQ6Ei1KhwR4qVaF2OZmaH0oAOc55pOn/nF5uhe
5+iZJ1mEd2X0LV0y3Td6ujch0rRwLauECTsLhCKWqIjry9D+mtW8TdaFJK4kPWDYAj5XFXj/7YfO
R4rRSHCCfhopMlMmFmlki11Q+bJIbhlWGryJ9y+DaBMKZSxW3CQ3TJj93cOe8BUkvmz3s3Hq+29a
i6vySKerevGvqw4H6K8EBPVRXBF1VzQonaQ4Y9bTGJJB1hr54Ecg7gQCkjfSrn9jv7RE3bgJIPNP
B+eQWijkkgnMC4b/w3Q3XAXP0BGdeS1axorYWMQFW+iDHKezsFFrx8Zu9ebN/hT/XxWT+Xgb33FZ
+lM7iLFbw1lMU5cIpzTuriPusvCV63vqhi/gTMjk9wMz08KnPLREbCCtXejWh4btxso6nQ0PZ2br
pIj2bZIXlNvRbFsxo0tWXC5lGJ7w5kTH0DrP7h4VUhWI2E3g1oWxnbT7r9dheYOyqk24/0M9rFgC
HEmO/K9ZCj2+/jWYeaGiarjwPaYBjquWYQLb6K6EbDwhGjzTe7i43tKZ5pHox4hzw+vOiULFglNi
zvJlbzId/gFes7Z9DE2HvOKaXMo06eDPybcFyoSWm9OWHpRJrIbNbbVFBCESsFiKT/Qii2JY9TK4
5t6TMxMA6G/w9WtRFV+3G1H5AkBs2bQf2dSL4zzNi8/IpuKm0jH4EbaSMobV8Zey6HLxNbX4582g
2JJeP6MWb5JY1TSyRsZqoX6d7RePxSa0dFyEXEtiXyAE3gecuufw4+zqxkL6FAUwb3kJkgSUFTds
wBMGHZxOHXaKcvQ1+PP9J14JAY/uw23Yc2QxyjHcGLQud6OirHkNoRzxlPSbUs01hUKbAZOQYxBt
u3z6ueib02XJ5HW4+uqgi401pMQ46vaPfB8rH6BQlz16xWOYfSTsYRXKpanuY14YKhmeJQMZpmCz
jOXpMxtwXmB/2wxcO95JDZFzYMTaCA04CK51dDRxTvoAzsDWG6fqlYiHlbJnvLfoTPT1ZRnzNVGt
DHvuNjxJ3P/MXtv+D6KV9vMRLMIxPb3Tzcps5CLq1BDDI9tBNYNQnqojuTGySN0AdmCrbSd//FZK
Rr20Ay6xjD4EzKgzWGgmDS/pIQeL/CFJv6iWxLE9jE9mJm4Nk6paJ5RhWhkC6aiXuuBeMN3MsJn3
D7+bzJ+kZ2jLFpa3rbS/3Y5EuZ8Z0rGjaBMGOZA4mlq7FAMmWjFMwPAT3riU9qhp4WRHe6tZ/5u7
4KKjg2INldukd7zE0KkrTQx3Z2nTvXBVStqaz4OTUs0Kx7k/ECjBU6+SD1ex0DR//2kdtGVoCHip
Do3gPavwGMAW2jCjCHSMw3yut3Id9fk1kqBsZHxa4X4UDH9ExH0ZH8Vacm02169Byljs4Cbq77Py
3o9ESgAtUYR8tuZ1mnyZOjpgtzbKlHZlvZImVczhHF5h2d/juJh96/ODZxgiObvGmi0fih+hKoYq
y2WTbynt6qR2TnF3nos0cC+nddrXx3xIGUfHXfTeMH/KJFDPeqgnwWmP5L36WzQrspJ4IiHrtiBQ
jUsYDay/jECMokLhshE2R1+GyXdlOe1zeHQyn7Ovh6LrJScySnY2GboVPkXPSrEGQeLF6/Mqav7Y
8HQ7i7LoSVeoWBk2ELlfQnWwlbp014kpNoDr4ET/+uSuEnzGxhfOVtZtBeL5ZU65knwxwwMdRb5y
LgN9OHBjov1rM9Znd+Jdvw/EbH/pNZokjRPDFGFMdZO1FdslxRA54YLHTmdPJ1sBeOAwfJQ+HCXB
Iq1ilh4UDDXCl1/A6yk758fHwqU3FJYHOGlcDeqjOMXB6A4ooqKkmer4EX8Z6nsPd5glXa7r21yJ
aBdssSHvG4DGEGLx4AN4P5MYVnTal2v0+vgtxdPie7F/CGng1jM1DPTdXDWP8MiBBlXaOqbWHbCZ
WFwzdwn/IxsdLnDQWWRg58NU+fSTvVK37BqNfTXHsTOLX8ntkPabM00Ir8zLXXdbgra33Xpa4y0E
EheuF39sm1Q0LGUhslPc2C5BOQryPTVbLPc6xESgyeTBaVBBnrq26HYFnDpSHVumIy9R1R+cAEh3
Clr/KjcftQL5AI9wDK9tcnRyJZqFNPlNcZB9cTB0h3V91cpZmGh9J9/vu5TwEmaWaXb/r+/kUZe7
G7T1r9hyA/8N36VvVSME8509wdvs6pnADw7sZushnmxcpUy5R2my5Vjc4V+4Ek6Y1CK05g/oqT6Z
cGWAdX9iwpm5aoFlbavsdGIT0xQCDTQzIWyFRviIxxV4Thd2bR9xcR0TDIVV7jEluGLxE1/ZwpqW
PI0tPK03Zg9WTkcpqylzpS4dxOEkDV4QNKNLyn7MXVdrnbyrvS0dPryzwoXiK+U9122BMARSAqlO
ZwRdERKlQgjozyG441iuQB0Kmpqg8D/YZR2gr8hGcC6RTQa+L5z65bie6QH0BDExx9FQ/GlyFllK
92DeSylYnhx24rwsWed5n+vn4LFgz6eD6kcmjsc6LWsyk7Djyqck8TtmtVAy7/izQ/EdNy53G01W
4tqKtZWtZLXwc3pPlynzK+Ssl6kAOysA8mbcyCokVVMGm0scgvjUBQicSrFSqcjHoFX4vNw0zFl0
N6Gyrj6vHIXiC1Gui7/cYPl8zLNDhEBSuQUqEoKybVbGAE/LHdS5Df/Q+kDxHajc/buY2mxSHtVF
GeM1XXEiLNh/fhP5I/yiV4pllC3DG4StnQQOkZAO2Uowc5K4m0rXRK2ej1NvdHGMqafx80X/iqDj
Wkkv8xONnalEfbMyvZDqMVHs8nRn0aPjtwEu2yNQbsiPlXE5MEzIB0GjMQfR9P4sb6m2NwCDM4tD
Rzn+CkQfe7IeRo2I5jWHE/+vTfWEKRMGPd3g3cfRug6Vmfj/6svi66A2l3BH2ijs7FfWmWtyJNN6
rKzf6uH/JZRXlVveN6uDPJ5T8xfg2xVaXTKSPRw7uvtuebvIWGBJUn0yF5/51qPVBnKFEQlD2KrR
ckrqqRxn7We7sQTwZIlQyxrHd9AQsQPUWvBXsvwaV9dr62Utyms/79ygkW5rQd6gtwDGqhnMfXL6
BUOfCnuncnNOdegpaob1famUbGClsOHs5543HhkU2crUiY5gLPJ32aWvaKipEmFweotK1jsrAOmu
jVdB4H3fmkaqB3J6wKsy0xjxEJ9uJVbJTEDelIGV0ugQ7GYkUyO4J7EDrZbrGifpVVAVDDIOy/S1
C0qK+wKrd0s6Mn4ezU3D8qqvaI2MnChJ+gDpfYrV2rgS5xHwCe60mAwUD7WLijAGg0BIRfVNBWAL
ipcsNXj/uye5NpfcguyC3be0dL9HDYpxjWyiJdiki+zg+3A0XjUwTLSLX8ZR/xn00bzYEXxaJM7b
lq+QzBM3zjx71r9ORRP2PMoOzG2Qm/0wjLbfkl1zPzeIyAWIEwWtRmG2o69yJ18IuwCx+/5EoBZI
MtvmGAYeYQcLoZ8/IdFl6bX2fZDZD9E88prnW3ccCAOm0VqYhv6XnlhgYZ1y+xA+YyimO/AHBhNL
IsF6oE4CT4UMMU6WpYEIKO/d+3tGjX9deGlnnUFZvMsdTNdBCw4y4j60R3xlJXc0I+Tg1gpQIyZP
8SdtF6u4ghZ+EHlfqPfej7L8c+xdaqDOzcnrBM5H48yTyMlhh7kuY4zDALeiZy5AUyOaQL6si3DO
DkKn8igPCr6CBpl+fm5AOwDGWvp/6NFAcBjkFcmF/KBThcyV4R+6eeqxWshCUldJP9D44+CxSgKY
ctYHvlh6EReaqv9o5BCOZ70reRmRoQUicQgYyfV4MY9YJ7MvZWnwRaj6a5iRgAwTSA+AjTaxzTT+
pJHhCvsnoxSHiVNuiQXI47oiennMXu+oYjNvwb05pJ2/G5nGdLQIDkEI0okxL2iwW6eCtMJtc3UN
RSxM1MLxZGhFxlAd52RyAGqp9LctYNwFQe9qvRHgc4eZZHFaFHcwt29YWZ/l5ilnPVetxFAn7XRx
iwTVG+vECFc/ldx0OPZgrh3ebcShFSod2s717ywpBtDyfucLFzXPFFg1J6NI30MBQXNs/RrdB5+b
qpM/Wmj2ofUoZWh5Zx46UbPpmPF38QCnLcgHtISN/CzM/vhOCCMLqGD3h6Qy9UfXaHXhDU5GabOM
4pbgPa3XX+CY/caW2dFb7Urc82q/iDud+g0aZlmdvjo/WuYJm6p/Xjp+5INs7wrlwNhycscSpsUa
PEmHanPk7GAVDaS3LlTQH69BqHBQntcQlhE04T3WDwhg6xgfTr90S07aytej19bv3q8cso8V6Q5G
L1A2OBTpftE8YqfO/wYBkPlcX+kyy/sSw+jcP9nxwHUtVwbgY/9nyFqlJCsKv4WZGvl3VysEbiZN
QMOZgppkJ05jsF3y8ZQ0fbyJMFtKiC2wzr5h5PM6x6/VduTAn+38Dlpsd04jp6T83thV+4ZKm2DP
4SjQcuCGIG6qWXxFCCaa+HJ4iqnu7en45/MqusSDCrMb+Fprxo/CERWsnU/BsVmqFYcqpeKZAQYl
HNEr5S31Q0OvHznXfHmDEVHRkZWyIUh0CAXeWbJ1vNMXY4ZWfsPam9XcGqFL3tUdcofRgAP5nw7K
riEE3Q5PZ8ZcrVK5e1i/ZpG8vfBkcGwNIxw2TjsVbnas8pQLWkPEi/1ChYYm4Lgn97NATwUS4jhB
cynpwuOYf/AXMutxk0ybxVvsHvfJbVXs92DFUBgceO93U13KmOv9hPtbQ6T3kA81MAHgehJRmb6M
Q9hLubUdNLeoNriq/1PxXPgW01ZivFHa2bG4e/loxKKZN5AQswS5VpoLjHJhUqK1FGkagsboc6i2
taEldqqQDfEwkqlQul19ApjMeJnyEAn3KJ3wKI3dxWzPFaIA+yEymPHUt4dSQfTD17xBh1z5nPQX
/3IrHNQP84UE3gDCPaZICyCgtbKbznlU7zi1PeUbx23JM6Tok4JgmNubq7RZHRRW//rMJ02cutQ7
yLRAJUPX5WUBh282XCZs7duW+Z0MGu7cOUbB2sIEN/uFpFCRXRJjUMpuRffKYm/f9xsSmw6asJc8
HuGtYjBEKvYChzpSJG6pDl9ONB7vcseuisR+Kel087DNiVFGxSQgWtDm19il9d1ufu6iHkDjtioQ
FaDX0xynhsq3RXcKowd8VfZsfP1G9FA4ZMCFEvL3nG85zGFUiKQVek82WVy9NSGkWsl/8D0mioIk
d1X4OMJNPWNuvwkkXzRtoWjV9khIQdQGnEe5fxGmRifKFjyZbq6yl18GHFUFLOl830QVgucw48QW
CLkriXl1cgEf6mMXk0OFpJj+hIi1vAd1obCsWBZaVwii40sL/TlvdIww/+hbLyz5cBuFBmuVdSlA
B3Rt1cjHDCruERyZ6B39krYXtrdX99LKa963J58PCweiVUTjpvk6J+DAEB7jhqBCGzmbeuAuc9H3
XqLmXz4c0KuoZ7247EC6LPc1LV4z7rBEva+lOinI26k4OFsvuiLx9b1E8FFx3T0NWQlCck0WoVvV
uALEOM0yDdSrmv1wEyVfWHEjhyWnDLMlYKWbvN56lSE69Y6kTa1QmLqueY3vbOMhR2ah2f8oeP4l
Vj8ugv88NaUIPBAxMcRmg0IJD7H3zteqUVw98pk9SLEUHwJXOB4/kRpNlt3KH7PmhmdPMpW85+XV
r6peaudG96+u97X+ZQi1ltvLxiryfJR4z1bCDrbJBLaZ2he8yzgSDJ6WtWhQsSw1g3O0sJYm/wdv
QiE0d4Y5wiX5jtSFpePauIKa698ELKGfHGfwwghFJJXWHBSx1Wd9E0thhmP9bK/Tvm0eBaaTvqju
12bkEnA/+In8i7XKyoLAllt7RwaJiOx4tZOfGnsOzb6i7M49et0kTZeXqh7NffUELn2zbIOu/33/
Ovxwa5uYHSj6lgJypLjvI4CGlfRbIFqHjuAcwXZcV0QvVv6X/Cmm4aZTdOOdPhBKpEVscPSEVsYm
iVa8gjq7bWoNftPagRTr+dv4Q+9XVeh++n9iP/DGOucoxnXnItlxD6sNPp0VzrLmNaTGT/xh/xop
/10JNUe9nU58lT5QUSYsEIGQiNgMmqrhxi5OnPiTCVoadvNhu56HP1U8NihYaR1lCSxUPWvpvWM/
8HPL40kPM3FYlHBqoSPDpvjksr95ZhTWbTcBYOJmbBcyjqUMgHG8SJzJeNDZLK5ZqxMrr9nuLZbU
QgR8BZ7WMgHdeO75+y9u6pCwmbkZ+AMUMym1oO0gDqk2sOpybFy+P71JZUVns0cnlA0A2H/quSEo
jwUNQFtZs4KyCgfJoYWEM48mBMcsHk+Mm6tFoY92lhYPSpnq7tKf2x08hJ4XiEOMxijm0/ukJdiZ
lLLtu9kTxKW4xMp50ATAJ5mTYmKEp9X4vlpv1q949JGwS/64HtZ0YCECxV4+MdVUFMKkOTeqPsZ0
GNcnWcZs/HSSPs2xkYdJqDnLlZtJHhOODHiPoCDiu8Du+juiJ8sWOmLe3Xval88FLVyRrDxC00mP
UegMd5Y4A4Eq2n8vUZ+SzyJ2trL6JgVDPg72n08BsejisphFAC4RDraIipMGk3FPK3/rxeo+i6w+
FXyE1koIaK5bLRaE7hAxeCAFpOe9fl/+O+fpvOYwxiTJ55AxnMYUjFQT/+NlM9Tg/R6Q5ZqIQUvU
V+3pK5YkcFmXQGUy17B5FcTeJXzzJ1YxBMARuonE/5AVv+GzsSu2iA7VFQSDykEbJIS6xV+dOE4M
6xa4n5EgLPdBETXgAFlHxumDw65nHerJwYZI1nb5p1mLGZFC5xbraMW/0XeCQ+RgnAc/qTJ7nZHM
qMAZeElJ5V+gw2GjzhZEl/U07WOtpRMtazpDTKhf1TDJeN8VOHRk6plROCHyVFDq6Czebc1Y3y1X
1dXtpGGVDb46M+si25vobTrSBbK+/5bljzhTNQAPySGj1Ie+w1GlZ3f0+77LyGVkRgmoOjYL6ykm
5uYGqR3owFcVPUzVVeopsMjbEX6mN7TyKgbZekL4OHeTxHuEWu92WHzryHPJ7YKbwTkU4ShLv5zt
G0p4CorRFdpkKyK2qZEEUvnh8riF1HUt3tRaeodrglgzpqKC+bZJdIwcu54Nrj9DHU61nykipu7P
95+s3tMc1bS6EpseGELcDIzppmAosW0GU6cGiaOhagMFTGC3W6kwvICnR5x2nmo1qTsPotJ6eG4p
8r798e4acmAx5ilbbCG/qAtF/9feCg+UEUjmWWVfgUHBcxpa7nMfMBAg0/WPGIFCdfggxF/zd3Qi
xOohR39M0DhebrjKbzrA8GWCCST9c/i8EHBFC1aOgoBrPtYyB1zelaxevFUkoz7AMd0FQTXstKwQ
qNU6/9irQ5MnbqVq+5rcCZ4pN4CSz9pIPvedJtiBLHQ2adH745tJex84XlLD5LcmnVWbMfHc0rvs
lYUCWOKMBXvs4BY/d7kK4SPD+kSdi3RfJgwntcf9Dxdc2mroZsw7WmV2N7qi6OUK1mTsoayH3Nzg
RzVo3crPEL79ezFQte+ZwApzLMrcG6wD7MdA5gshZpuQWXFAsDwSkgshFyabFyMLDworK+rZZm6C
JnJQ2g3HV2rH2s5hLpJZ0vLmrh1lzYS6qdnE0APb48v+WXBN7w7hU8eu7zzzjj+72Myfy/1W49Va
8Cj2LCH6IWaC3XDNIr9CX/AMGRfEHgGguwTD5azTtv+QR0WFzIU7NgHjIm1jj+Eew79aKwQu9+AG
58+9lCC0/nN9tUByhPZLiR9dsj3dB8pHYJc7lUiKJuiJFC8Kc3M6CfljbQFguHNYkBlF6/GXrHGA
s7h+ZaWELfnkwkL5vPIg5vEzRK/xMYRnqfzCgxhNI/3c3IWhimRK5/jQeFaaRWqbSib34yO6p5qe
WlCDs/HGXOlyT55/2j4V4hMCIqCp4ARrI3SJug1JBBY6CkbaY4ebE6vwr9G1dm5V5/Tw8iG2w451
QipaX2RJWWdLzW60OZiMqGtyvxv9ybxViJCBf6AIXBEuYMQVZ+GWrzVJi0KkQ4M8Itvtha5lbyWl
3lfjM6jrXlf+07mZsk/NZIWvRRX6WhTpA/D7SD3gB8e4KfW5iuN9vFH6/Yulkpp0Bg5vs1je31Q/
bNhLc43P5k67gQOEt+Rhnd2GrN2ACqVjozIGbdglsVYY7LBuFTBRyiX+lKoVIGdzlW8sc2p16puH
aft5S6z0TBa2KuRo4FUs56rkQKhUdQY/t6V2Zd2mKdEXN6jcslcoIMFFWkEZp9ZlEOrblj3mxcwZ
81wyH59xrg+XHzvLjQDXYJp7gweVjd2FFIflIOqIB0JS3gOwlhm1WSLVHos3AfY+dcOxNoTOHbhE
+i5d9wv7SR/G29K1r8l0ETWq9fmY20E9+KIuY7hkhyrfaReEHe/8slc8U7PyFlPz33GgMMU/Ibvg
fm1HEdipVJTCfTZJI9kXCaCYq1vmN7wapKC7VmKdyRzF96x2+tsBEdwv4QsaNNZHtmKoBr+ST0fd
Uq3MC6rppOFwNKPxTIbqfjG/ZLZwApJInbZc3z+nUyuxAVzOslzIWOHRg8RLcOIN4gO67V7uZiO9
sBMYQJ2vuWTU3ZK6wdt0fpB/lT0I+gFqzl4azmZtkF/9hjvDPtYSp4o48gJlkVg1M7vtLvzkKEAJ
9Zz4IVEWRH982sNGkmJW6IYUuj2p7PHu3qdJZp275YOqYWPTkty/WAdcJSB3wvV830XWOVfD2OoF
NY9YVNSIP/dJoDBfG1lPALLvEar8lEG9mhcqPplWsSnXlH8r660JEeRk/4NR/MkrZQJs9/ZBpLmD
godVpbXfoP9EO16SmaiEa7nvA9nJcd46hv1ame/1QgqC0MGGVLftE8isZoH0nlhF7L+aGNcm7t0f
3LHoxqeybcjzDULMdYvHyXUBOknUuWWBpIzgJ5v9WilFQsngc9UEVfpB3/ZYSeVR1LBbajONhKwQ
IkGYB4QB/1t/zyOscDfgyN7XFoo+eKH+aLbWpLs8HzHkbrnJdSgmrB8GmvyjdgnBKSNVpfRe+4Ck
kWoGIhd/mHDZBj8SyU8sphl+somBJf7NkQdV1SHlkWsnWSpr1HKRutmxthopdEvudDhwA4kI3mxQ
n6FLDsf2UyKNHfDNWs1/3FRT7nvmOEPz4HEx72yccObzTLR3J2o5RIxWzUZbcknrTEBSg6HNXBD5
pSyQq5ba4UvkFZvNg57WKE3upMbgntVQVLVTUrug7O3ekvk/ZbpSzZ5C+a+xAj2vHCIS4RfsfiHb
9ztFaAgHYPyn3Uf1CcX26v4cFI2zjGZk6WHGtAYzutw4IabDFBx8339gMMujHsg8dUw5x2+k6wXZ
185ozZ7nDg3JN/idt6eQ7P52Sy32FEnTZgItSPG9JP3Y2VwawvCmtdf1ZxMfD3zmIcCW+VXDKyfI
vZJZEz69rqC+7I7uMDl0WJy3o5I0G4pZ4scnRnslcdzOWZHvzMXpHRzNOIB2C+iEYlt5iuc5qoE0
w/folrDtNHJKK+CW/0pGu7gDXLNp0ds60U7oLWMRJuXiHReoeQF6OkC4WfEiG1OQs3KvQYYv9ijx
FdtkdkkUKjsNv997Rc8kzsOKzekazxVBlOuYOtWtDyrjLZUtc9UbfMPLIXlCAd97vrCoFEch72fv
yX1f6sy3WNmvC8v4f4px+AwzzIi3ULFEWAY2T5/Mx4fZ75f3T6VpsS1lc+e9wPN7iSvXsz8c95QN
B6cAguMrbIYQ6ubQt3iVR06TrPQJLALnmQpNSqyXQG8a9EW20aJnznD4X6jrMrGuhaAwOEzb05gi
XVUOhxpHLPhcbUSKFGkOiE9mUjmtrsyBOo0nJbq3p3mmcXULBJdlouOuFHoXuw9bE/KUyTNODjHf
c+fXgoaq/nwYZE8qe5V8ySaJFYDQQc9Xn6Zy30Mf+A88kQRq1c/yodY1BHg7JL8BbgKwL6aiYEB8
RDj1c7i1KnhGm7fDNvLPLiLPgww6SOYwHcbcinBRNU/frv0RXnpIT+JMRgmgAL/bjudTsXT/ibuh
ZMdjbPTHWTSKex1aYM1LzSWhYtX1JfBR4Rv4YWjQQ32MbAX0E+DSM54U1B/dBnXrs3kKdHKjB7zU
Zmmi+SGXIDWWFKGiZMkbqX4q0Ift5RIS2sgN+IlARAb6cMBOJ/+vVJmOevFi5ZmmTw9vm3DAHz6y
yfLL2hAZ8luTQQkZ5QiPFThOIy1G3yMBGPUzMUdxj0l3Ti3WVywMlnG2tfHSOkedK606exCH7GLk
QvngFDY0OSKl7bE8ho3zbDz21OdwtiWqAhZjrxW0kWEWbbnzNX7Bd7qU5+rvxnBHRhNN9FTLhOQ+
XwvvnYu6mJgiNMLJX+1xJKcTDn5QO+y58T4T8u7FiPi4Lj3RuMKQMUEzEYrFzMxPfsJIo4HuLV0O
mZg/MyAiuerj2CNSk3WKhL+KcaouJCcI1aqHZxu3OCI9pLaKp1rsvjY0QilxX+ZrBf1Tkaqeb03d
iy4Mw6uP4eM+3X6ghvMHHDCKXrNKCR4ZmI7R5PBI8TpOFuGKEz+axrQooSHIvHnx9TeTN1bn/FLA
dgWjUqFNICUEyxm6xdYaNzbpH+kh3yeRWYD3xGV+rVkF4SDCnK3BELMUlBIm5KObl7qjww6yFXgV
U4Enwcd/Hm2qWJYxkAE7DZcE1hhrdceoY4NFFsqurg0K/mHfTykbDx2Y2ulQK590C49CYj+440O8
11y5NCf4/9tkHCGPRErrM00Rr+oQIgqGQrPJXvOTq1WmUHY6ikHXQ7tddBNoIIIhRg+Lcymlks8l
fAFNspvazwUSV+33NjF/IQNhOfjfrVjRYNE2wFt18Iy3bzVQ8c7n+wridyoDIBOkkM3koiBgOhav
ZtWj6gosTbu2sHeAdYlt7vNPA21+3M74+aXJrjxhjVgP0gf1NyFXMrMASApYCDoOQF39pGgyJbce
AOD054YZZzV5rVIkjFmNykScVQO461j/7De4up3JkPljm0cAJda+AodGEbcPhsPIS5y2wBZgqIM4
yE85Dcw2GzW286F7+aBGOC0rZoCOHJFS97gnUONuEi23V4jHTCpvD4ilaJIUf/ZNy+ujVFQYdskB
ewu1OT7x9YoUxHF26+wCh51T4JgzSriFBP8llpigTAn+ILgMxAIUh3B7SzB2JpXAzhYNLHvq/kl4
RUd3KE/ZPhvLlihB6uvB6KpO08x1qjwpipbeT1g+i7tIVdDl8z5Bfcj5Av+gfrOogkYsNVhKO4pX
GivJQ2zWIKiztvSvgzT+Rn+7XY19bhyy+oHbmoYOM3ZUOoDRmgOg5mH6OkzjWkagvm7+IOanmH4R
/L4JwAI55BS45JHf01WT/HYfGw+7l2LoJ46X3IF6LO0EK9+kEca+Gl2x5RwNELJdUTHsP1EkjEbC
bMqtMnddFDsJBMfzp08/EMmv1ZAGhnZF5W6y1WdwkLGCKPu8/Cqb0FMcteg5XmMBhCWGoHQ/t/5Y
ZQ/nkYCBEf35LZTHtj1KZc5/7YqTj9nAnpOiTZt6Ed9H03ILqEduXmH1nMNA6HBuuzmuK4+9Xw3N
hVEm4I6L6XJMO0Ap6Heki+LlaCun+lvqxaP2vNa7IyzqZ7QFAwanF7lRzbcz1Khu6q2+UJUPXrnT
D4W6+4HFRDl7Z0z5CMwRkW9GvJYb2Jzw+f1116zcz1Inp65DlOJ8mpWuAUUvbDkl5KNqy67rmKgF
F3478PvdoZNxAaZceBXgTf7AGwAxsxMlkEp/BccbwAXiNGEPxMpZxUM8ts9LgIcti+ZD04UmbPno
4tWCv3QMZwE3RTp3Tf7PnYVV9joQhDS6hlFDt6SfffyrdhARWAZl+2fUuwZkIaCpZaL/JZ9qGcUc
9+zvz1RpQ4ef8wYR0uCdYH8GjCb2qQut4Ok+NFQykXl2Er8CbmWPWsjwkWYRC7IITVte4aElXLT2
0pYvG0GNKTRCr1pm/7dfS0ogRJI89g9FAMG0FBZo6M48ARPYbwkiDeETsXgwfOW8POYtMnny+2o3
ZHLbxcdzgu7kTZpxrdQYmC82Vjzal/xL4GcbU7j0KwFsD2NW6u0rzeR1WnWA8ZD4ywuykp0xau6B
9hW6KnizsPHIVwPS2HGSQ34w+i4Yt3l550Jwl6HZ6aH0f0X6TkHltRuoSKkxIv7eDAeIlBs6+GH6
93CwK6vcj2C1w3YAVIcHrl1+yCIZB+BhUpJtyQZqvm8sDkMfJIn4HaQP2Z57GzsthZrL21ydpGMf
q2py6xJ9CWqkjeEKnE5a3XexT7/ebf7G6EjPvfjN6SzMVtj82FCfZKMJgodCE84wcUKcfXLp6znD
fgFavds+0KISle6E3QsQ1RWr/mFGEcFNNMO1af6/LKvKD+0KgXKX6uhad8h7EGIuVxuEwWfw2lE4
TpryUc3P5PQiwSlu2MCP6Pe1swPf0nyv4fHLWFNIvmhdXlnrnUz1QKJpsF+vEHOpQFY+HmIJsJdD
pUetIoTaVoiT9WIxRGYYjQ7MV9Rs8CS6EanAMLIvg7eBGfVw22WSEJpHAv0wK7vIJhiSmKjG2jc4
KVNfPJql8Ll/g1fRppsySZsER6sxCV4R2qqZxALDD//K+9Xkcu0yWLj1vN9MG0669FX51eTqRs2U
698RL6xZH2KQliPxY9h+9eYMztyH39sBuIOgBJSNXz7sk7BMvxsDNLjp9v+DQBjNMX1Lwa7T55c8
Rzu0+lDuSz0FAkBCyzbnDJKe/Ii4QfTMFsKz3Q8uemAflzqlhMUdN//TakmS5TYHAVn/dqUZw+fl
2f3DCLvdFtIYnvsss0RZm34QwKySZCcD41SvuRO3/enY2zm/uqbwCG1wRrMBuFyIZb/adAmrmmdW
CGS4hl1bQLv5jn80fF6RftV0oU1ETj1w1oPYzVQwN0ZUF+Hzc/HLf1AWsIWyukPLG8CwOC2j8Reu
qpsd2hSzuHmq0U2F8ePClniy+WwSIGGXS9qjvRo3EMc3vyKiT/d0YQOCYZK/VjqtFG3iSvFef2/r
fVOfn/g3+UT2s3OfjSq+MfT1Oix0zSJZX9BVcs3u4apFit/UamOtJCo14BTWeo+VnjdQnZoWdwg6
0aJRiOiFUt6+7IXAS/GVz6SP+DCT7Z14xgQ98b35e/CIIFi6ioiltH0ZifwkhCWdsO0iVvTmAHQS
OsV3WLWvxUdxAzd/S6Iic53dIUxWk7hu9srJMZqYw7qOflEEusrHKt/NbelB4tzOIumkjrelXpKy
jTCsKMMbZZvA+vup8vlaIFKhv97TuHN1McLhlgAEDHAk/TusFWmTwFSQS0/O1Nvms4W0COCzp7P6
jI8mKzSgdoIBlAPOOQasE8dIEfgMMRsXGnLr5WZy20XDyx5lxxmWjvEYW8Km/eYGFMqlBCI7gtMs
M/fUoYXINCgNGwhwpFR6IA3kQLN08TEsh7NligUAaNNn3jKwjXY16TK0rIoHWw+lhCbI8R0JtIfM
qcWgIeoK7VxA8DiUUULNn+bMUC8SvTCuCI392XOOxnkD0GjTYQ04CtDil/aU5BFij0/s34FFw4Fs
PQIIxUJ9bD19cC1n2oIzm5DkwyBAe9uSTkGdGVNPa0olZNzM1WBNsHrEv7GImCS9YO2s2plWnKnX
JBksRp5HlYKpR8JtDNPDprnw32xyhYcRc0eWtXitctp4YDhdaVOv0lKL9ADdT869fvfyh32YQbzT
qWrK/hsn3f/B3amfH+JOsT+PuOmC9g05BPPUm4CkyqU7eY6WNFtVjf/jd3qoI1AuziKGfMAVF9f/
SvROv9eSlJlSFAYaG0ifkjGh6eBFtBilVcMWpmJYFbEUAprOYt2BopZA2uTfFshWTbvp65ZjrhEx
3o5FmLYUnEAnDBPNax8cp+O7vUYAgAyIoxSCi31a1tvNRgd660dncCk44/SNOxKz78bIzVAwrUb4
+pCOY41jHICjmutF0CPUsN1Zv+UUdUmXZ5UkYGdGRq0+LDaQoWsHaZxFz26+4Orp37kCvR+Ia900
WY/fvIqYLQcJIssNMI0gXNv5BC6T7fAgPYyeYa2bOCcLbGVZguku3lboJa7a2FErY2ksexoHBUg1
aJ0oOLPub7CBC5kVAY+nE7QZu1HXfqi5ZxGWfcO6XggvQFsNjMOozSGuU//bxPDOZpsFyDmNcWvd
tfVqMfOUHcMsuoaavEoSI25pQG1WtZFlF7P4cMXlu9k1MGeKRxR/zKN5KEYo/oPeoiF3FfuFrmEA
EBcLjIqwXyVqaMmrLD3aCkk8LhZlXE+y5HFJBhjXH0IRaNwK/Vp6/5cH9HUvyidKe53PhTgR3mwI
Vjb6nf+Q8ByLNBCHA4fR5NUVFEhuGhZAdCsNDsT95EVLqQfpMob8IkMrHZGH1lagLEGPuGhZnLTX
w3LFmx4cV3Ddm6PVJsIEoR9XA/35UcIlc32SsufkhcMyWWOP4wkPSdL4Neq+8K3W0UC/ssHqAt5F
zg1+DsjmBdH4i3PVdjOQ+1lEn+kpp/BsR3fuibCeXlqS236n6u0wJtbKr4e9knO73ErTG7TkCe2r
IuzZmqfG4Y5MjxmaBGGbyha6pnvZAmVrK2P9at6tHeVs08IDqmQEdSY/UxbctaMT+zeHCFT5X2UF
v5VEiRywv1v95wof7L0xFrkV61SeRbvaQ6MfJtRMTISE99nvV4HzuniauiiFhEEbXletpm98ApAV
d+yrBNbDgasvCMuuG3fzLsrHuxNJ0f53n4aFNWMuYFqlwHFHvK355Nd8p3D2ClZCWnqi01ppTPry
DjGPxfrcOlaDnBgbME30gzhyLzzUZTe/e9yHpmSXLDJJjEbmDSsYWhiW7uHKWhFrxH8jBvAebP7u
9V6utLuXmeiDxV0RaTjHrSZmar2ruFBaZ6+EVoOUU391W3sZvmtIif5XtkQnLwPQmWxMqkvarOgC
qEPElT997RgRI6CdTCTH7hZzqUZHg+U961OVgT8M8Ty6sk6wVpD9ShtQR4mkHlmRqTf2nPMu5UBB
TFasYCW8jD7Yo901s6BEYXGZeibMAYJPDlLJd2r9x6Ukx0qCt6eReFYC/m95pVl+yGegKvsnbukn
OK5Auf7UYa5NFtou4s4Y2+OXmAS8zJJlpeesvIQTHfs3uR4tKg5BiyPWGgrlLYmhN5g2iu2fBg3H
+IlzczdJHF+UHTZupTf3puYKegGAwGYJ45FRN/c6b4Ya63znOcJwFNQ1YSdq4CYTdZ3wh6iQOQHZ
NyyaQOJj3M7epfGtARTBfmIRtxDTpgxWH+2mA1JPaMJIghFujzvEZ95kBupwz5pnXTiKKvV1kDVn
VUi1CRCgswKFpw3IPY9OwrAeq5QnmCvznNEo8uLY4z0iYl87Wdo0MZoff3/Yy26hBVsud8MwpTm6
k+Go/WUTRTGpfCWfiQSPrC0c0ryWXgZ077zs9zw1o6tH7UQX5ddvFgcimLL45Q8WYhNjyIZw0p9t
Xg4j2aauQAEyAxWiCN7y/2Q+/wbNBodqbcHSS4BnnqC39NpXJbJaiPX1oNwS5jc2p+O2GtXS5zhe
Tq2oYml0BTpDeupqpKt24HKsERA8/20gwkfJIiRaCWUQIVQYgJJfsdEGij4KuuewmW7pmmnHqs7C
pDjVRum0qqV9PPm0PKhBYJrbYhE2Xm53UWcaOz6RT77dY5lp+DnHRCudKaulHKhYLwknColW5Lw6
/dJbIzo/viPfDU3+SUc59WCGhvLPSno4/pKlPATrcWUK7+fJXiZqXat9y0IBu6ejvnMgXhGF9RRG
7P3htwTjOk9lFhf5pLHvNaelyxhhexLmLn1ZJNFAtj8LjneMBruHIvWU6cLQTPP+ADnOVF8poJfx
ZT84ANQqanEo/uMC+KgCJl/l8wfjV7HT6iOeNJ7rnk0eF8BZWhgs68SA4TfVrRkkhKvdM/9uGn6Z
/VsEUOlEeCXSGQFO4bKWeVnYo+66GfxPY5iKS4elNco1J+zkWh2JBdjT2MBKm5Zlv0Yz+OMvwI5S
rlRf3UK4qq5A8gIvYaZ8KW3GZxdbXm7kIyaUnNcay552PX2etQgStXEsdKl1NqJrQApXnm074UwI
QCwvGkdEDcmUkOGFK6c+fwlyGwGQ3KsA8epDqjKju1qR2O1VH0QVcD8eFHOwdXSCAbi64TVaci89
VKaqgDsk3ssbBGn/0Bm+tbo4KFwL6ZzeWruI6inZCvnFGwei9ar+pUyZw6tfXoyW6fXZRMpNDQ5t
nihL2PRkB8RaMHRU1D9foiWyZ/UooNlxXLW8loukdThT7Nr/8qm8aBTxS8hDBcVcMAtZsgWoBQu6
BOn854FhfcF05IpAsbruMJptLBw6VQBz1d3+WK8xeq1iW3f1A+XmwfC7owlyBE0sEEd4cFjDTUMb
tXWZDEtwXEoGqPc+p6JxHmcgHfihA4OibT51936jnbMIxW0klxcjnZiOg+6iK1RY/saXwnpII8he
rA7lGFI3VnuHO3w9iTNDMXZRf2EivrIP8hv3QppzVMA5jCEqix5qaiPJRn3A0iJJseAK/RkQ+2pl
B/Cf45lj02ydgYi0L52RxZcezolZPquElme8MwRWrGwYmwTuc8DwPmd1Cm/8HTddmcNez2blmq6c
N0dcdIJSSd1GRMmHbDH2eqnOvSELhRFV0zqy+tq/W1KgR/+xLteeUIOcB+NOcMTfk9UopRCob48h
vfOWhqucf5aZeSHYRd7qYnuZ5iehmXnZgQuo2tWHC6hupAMJpzlexOC8noJ47ewd19BME9x4MkBS
ym2+4C51pjYU72l2sPvAVe5UdMy8aUpRuvTrSmUy0g2+Qc6sbvJ7WQZmZDTDSX5MHyi7tZ/dNGHs
8uVhOgIpC+HfUxEydezHqURlT6VzrT9iXbguCWRi5lBqO4gkDZ4+Ev6gVogTTxo5HG7eCkDV/qq8
6C8doAnj9rA5utuqfLtg3a6YemfkCNoJU3/5Eq1tpw9ehySuAjlX0PdkPtZPAvpzMiwhmCswSLsQ
KrkRwuGbjh5FqflM1sTLSHBWSVRpWip1TlNh7QhnieWK23KMjVoMh5H4W3IydgogAMld1DSgL6hS
bX2dDq3/55n/yrK3j2B+T8b2hO7+9FpuQi8YEEkFNEAkAKMxaa1nxkxj6kZcZMO6gr6N98P251Ow
rgA3rlhn46VHSCdWZqvJ1pNGKK8rz/8q8+v3WcKEOoiKamj2613dI8fQbU782X1SA2pzZQ557Fah
YJqsUxvO1xFqYA57qK8YpEVqDCs+KqvBzCUUYdBwGDzn4JJPFoFIFgqfqU3RGsj2wco4nx4YHos6
sV/zi+6ek8hz5rdFctTybkv9YycFkY/Hl06t3v8ZciLIs0D6UzUI9miZhcbbiCm9ur2xr+TQxLT4
hjXfrsgUBKku1A5u9+QQRtsFAL0BWyX1igyPf8D/C+b7Bh1rbaC751IB6BbpGuI4EUQjTu1ALEnF
YbsM5di1qO6H4I7Yte0/5uTCRkYNcP8W69QS08yq1uHhW/aGSedZlRsRzw16uOABigqnyI/5Z0qS
eZkMqpF5nXnf5ZtUDuR22/KWtj5PY+jGVyTMb4/TiHavhmvgdtfzqq0dQ0JaW7vyf+RFZls3bVz9
fb+4VleAxmMa+QRvvHu7cNRwEbfC3ah1c4cFVr8j2t880l2eJsQ9ub9szdX9u3z2ZgLWP232nfTX
BacPdyrJ42/MAqULIjs+y9a+56KpVoTXfVkUNn5EzlizJi31u/5omiofjE4lBzKN4xkM7wykuuSg
SeUn52OjLs7aW6PZHQg6RiUwkt456EU5fynJdouhd0jUBKh1LVAT21FMVbBm1KqgboGwYEAxUpOU
Mevr5BRd1xJ9Rs+hwTMSEk6GCPnI2IxwecoNMZlJm5ky7zsgyYsvrNEId+hwATDZfIB2tp9Vz6fs
7eDfoidaAUaKRZy/u6ZC1zauvXj3MMdn8HIOzkPou7IiEMdeTMmjB5GSJi72EFbd/mdwzPTUPGws
YGJtPRVHI9T6apzWgFvdsoW8JbRa/kOQ/wzrzh1RL+hz7/kpgDgyE5YJh4laGaQUfHxRbkIlDiHm
UvCY0+vLOowfmTXU6SLM0NbaQ5vb3gukx0q9PxFtg4gFpQemqAtqw4xEKvt0LYwuJyiCSQZwXg+4
5WLkOviptzD1+D+o3VhP6t8sTBZXxr53/WsDKVuH19cFXvKU2eDJj0dP+0YVEjT5KEMO1EXFhG17
R5TWkfUuKpO7nBc8ZpB5eMhfL/A4DIQ0FRAZVC2XoKep1vEQPpO0t8JzMicCf8PZcsfwzWme1YcT
B6D94AhSKV7dMMX3Ce5g7ta69W5NNHS2d8+10oZDA1qaiR/WrJZG/+Sd6jtHtKtJqs6n5pDtqVWn
gXV33fG9vPnT3ksBnHIfKz7ve0WFTSZ6zusxXP4CH6gISopTNZxrmv0ykAzjctpGZa4eW8eLy4tN
FbS8lkbT+GvKFvdeq+aGijm1CUSrqdTESAQ5dFfoUDoKzCFET6cAiimoaGE696+t4Q7qmr1NmCUv
P2lbW5w3kddhnotqZAb9dkX7I1yNNyzO1E5iYRWvxiy27by4lnwaNcHFpSUGKiouCaWfBQShKJID
lCjYa1S+IrJ94V3PPoXUWl8WT1MHcUwCef3tqrpe6eXBMTmUboy/mw1OZ+zUUA/NfAs10MbAgzOY
B3B1NkMXK9yIa1se5SX3UmlD7RG3GhkgptfXQkPSsioNAsFgEHRCqOVrTNN6OxnDd5Qv5jjYRCyc
ObDxqUfiN3OwYEvc7rUSJ9HR9aPp373G4vYznPwTxWsvTL1hnBY5hU7h3xAYWSDqxltmAbc7s4e0
XZVev24UiLx5C1wGoVTl9y97FRr5t2l3q/j0/rT74ziWpDpxiFPdLHiCO+JGWm1Bi2TBptkibNoc
ta2CRpMNZc0Rc7QfhgrIEPAQo5TYGlps38OUtKovMlnUq+3J89xVWo9w3mHruOQgWeUywSkmMB5r
vaIK/k8IKGjrauFObnwuKT3vpY932ed8bRBxRX9lULJxBQ5L6jCwjOHiUf3l3lpUjC/oL0iI7mM+
lDcXoYAEThhkdSq9jIhSpAZtWrUeuFvGi0hcCdRfX0iR7oE3W0X0dN6moeNLoCcbRoP2GCDz2edR
EKw+KGdP587CfcE0pDnHPgWW6o7UfRXKOEh6HZYs61FIPRZMB/Mo5dj13XVZA204Uc3lEqSeu4Ff
PPxfCMCnLbHsxycdlooMlCIUQNJGzptdu20HUd5bqeGJWcT06RgTjJEJpGqHVC9uLmFW0oQrY1j4
6LasBrNVfkLHwKjGukMYYp9zFIJ9toEWes48NgolZZaLuNHqCXJLjjHMtx5H2DnNkGWoPYWi6lbJ
CMWJCVAtwI6teuIeN3gppPXoSg8VFigs9GiupjiwHI7JavamiyFrX6lAKC4q4ehvnyyfcsixSFpe
HmvzexRt/nKkXWzQmi83eyJhrfmzxIStwtl5WCqdbpAf0pc1oz+lm9oA6dj0WmwlqnurhxsX2F12
hqeSGYfC0OXrkzdajCcH3gjq7zKUSWEV0RntFoX+pelU+i7MzD3AEGpDUxcP0ymnEqOOJrv62S60
XhaM6/2WKYXYZMNzn3lmISvHEs5PQjZRV/SqB5EstqMrvSxnkpZsA6szO5Bhqrz+iQbJHQ/6Uz5g
Y+C1zaT/nCMUW9KQX6eymPUM7zHyGkRnbofWJQUH3JTAWL98nvSzC8LTr21Ck5759SRg9iUbL3+J
uvoWkJLgRscuFuwNXfiylo1GXKHjjFX7OdGcCVtZpoWiRgBhnlspV4KgP1a+MFKwzJgQncUF60Z+
mxYi/cX0nuRa6DgJt/xyVDuD3RvkRPKCf//xU33vOxd5tYKlXK1P/CwTL8Q6dlrxZBfijrjRL8YC
ncsMStawpM9+EMKt9x6U4R+/MZ/N9m44fdhNXCB6Yhoi9NT23g3KT4wnkV5Z8JV2PjWiLSq3yKC3
T0yWUiquMcc36CArAlmmLGcdv6vPOSVBuCzp7nCeOzCbwTP2xnQ+GdwjRcCQWsQhoSUVcL8ZYNT9
U/cwSMLJErKbF8H2zRzNVA0FmvkovHws1YLKPh4LCwnjyzBC+k3LToBvPFUPb1cjjrrHF67VRduy
urFdlFINVIcR7qILKj9nzJq1lodS3GINChPPMaZT/2XtsK8Yo6vHs5DjfkMlPL/9A+wtd5DtPdfi
wiY0TDqaghi4RZPTcXx63GRD7SO4C7IgrajDsdfG52l7mPhnwDybrBfq4xlEirMx1tKKx1arQgcW
BbN9If8GLm64aMUu4v40Sv6bJGLjeAuL0U5HYuZfVKz2rW19cagw8ylWL2j9WLWor4IXZtVefyFS
MpjLjdsZjTBZBojoyELNI6dDAiamWami1GYV9BpcNaGzl8bXqXnm1pqXWCvsg3UdAf3UKSHVKqr7
8GX+y4Ud6JCL1ykS1r6VgfMLNxVRB+7oesi3k67JVLRJ8zCcxMQVJ/NpVqZUz2wsvqeXTXwn+S8K
ada2ETlKQH7ARhw/NxVu9tYZbx3Jk0nSgiJOlmWLUG/KJZdsAiR/nb6B3sam8Sklx4aYDXu2ZuMK
Bb/SkP2+Cqag5YVkcfbhrDfGdYLzYi4VPimP7SFNjnu974xroSJVamZYr33Wbm3dqn+qxzh19b0o
7iQYTXWGu11OHWBB1icCTPtdhgZ1Z/kPAf9KiDawuOYfvuq2I+GrQ5LbsmCmG4Ta1EhC9sOnaHdY
+kr/x7V/o5kyYAR35rxTX2fIuWmrJ7utDxDjzbMtItpu555oyPdAjOj/voeli3IZ4vvqLYq5a23m
9Zrt9thDVwghAkBI/U4oVAkzRQnxe6N3PXCctRtggiecL/wfgEXvt03GtxYSfh/DyojCHz6OlhyU
yEzJrz5eTwkODUPIrZ9ECBPka76Va/Ql70AOnCJpZA68PNFVw1P5XvkA95mdPqu4I/QIqqAfW7S7
HtZDqL2F2B1H4Y/oJ5HAUkm9tpjNqnrAJ22e3vMUVWqLEwm0TF7ubCkH/o79D6vuIYdh5Zpuy97z
JVoep9ho6wy+mrFfInWG0uFSw1vawjpnNqqbIAejQHFRtWhg6gXYP/YWwHtmEXvdHMGLft7EX2lu
1ZBwDzX3i9wXq8DS9M8wgYE7DxYcXd3huM8UojAPXcRAdGm0L096V+jaso2Rf/9tCxd5m6Q+PiJy
afs7O7YU32fpTtdl+bx2UulB7Z1QP6nCugJq4wpFDXTrifoGP8mO9fQJDUyi30i1B14pUGQ/+uuk
+v5tTOdz8nptKGrZsCrgfQ5/LKUocnk7yIETlS02s/G7Qd6qPch8cpw/1MJfT128hSgnUOTVVHUj
nvAI0rIu1kGJ4SuCQutwCGfkYmgxN91ytlNNn7GIqyDSTL3wy1j+NVNSC1ELsrhPwuCQUVSrfd2b
uamUDxvRj5b5Fzl34J+XOVl1ZOcRAabA7HcztfcSQ2unLP+73CUUt3AsbvX3zhKypJCnLl5nkOaX
4gfR5SAdxj17wGkY2w5qcU4nKFFasmq0etQRpz1Ash07VTorTdULTutXF7CevvVYL+G6jGTCFvRL
JeHI2WUC0IcoIkKSQcsHXy6kdgy3KUwYr2PiHgwOX7psRZuFzKxNXUfopGjbTy7ZTlCdbizZKzYP
5sziUjH6u9+SV+tvSFXq+pSUClyto1IvANb8hpYfWh5c+BMN4U7SjkxnDq1v9QOqA8MC7QQnUTv+
jwuzwQxZ2ybZBV7bEi9G0ytBXLCr5EoLetLq9yMylGV2RAF8V5jlIh4wufFJvqitpMLhiqSeVPgM
rcL90cNB9LMiDHzmURy0F1lZZyuIITyFp+sohzM2Yz8ooySOF30C5w1/WlfKjWPyKfaH6bu/HnjW
A36tZgxSYAO2wR4PsA5cebAWa0/yhYJHxAFGtO1/9JlICTIGqc8ldfc3wtvTPgqdAViYBR09Ehgz
Ca9BpGZBquwciPJfZoWAqW/9tp8kGqxebHMLtl40AVl7tyc7DPg9rDjHHFB/KuU/mEIVMlk4dDAJ
wosY4PibDBv1A4WdVAuFJgrsE7y7Czy5zeZNRVe2so0aMLk3DD/CchKjr9fOXus3Y9KOm6aN2lu/
KkRlw+J1ZeE61JAI4upxzmvq60wtpCIboEV6WJ4pIZXJzk91/KQtVy0lcFl96QusPJ9tf0LYAxYy
n+nEK69YCyC2ew/vMl9VljtFcRoIShG1JZK1xfEqTfOV/y2uj6hWRXYGbCBEsmDGbMc6kdI9ze66
fO3/EE+L7q6DEOKMLF/+188Hu3BMUH+7UQhh+OKUGetdmZ8mlA/b/3Bbroc6AFLdUrWxj3AvjxhL
hFL+0Ff2S7nBEUmamxbIEsBw332iFVMnSHuvJGG/pX0OoOhLZJqw1B+cbKaK3JYiFvaa+KmPs5iG
2B2gO2u5/CMnp3FWfq8508u6Dmy1Bc18K0OX/aqj1I/JiZJd5jZvBqqztV0YES1wOxO54jEoAmq6
E+LwvojBfdM6mphF9VgYDfkLQj2me75rCc1RApIXbs7FF5Z1KH981nVt2sPaa3zsprt9bOxVUJ+w
IJ71cTP+xrXWqevCSEquvAhEHkyP6qvQZBJ4k2SZkklKqBeyp1wnXo9yGMwu+44C0g4n96EAz24a
39qfPY88ejhwpqAP/B9AEhmqxEth+RWehFI5htooZ0lwWGGGSkRTM6B1i9BevgkjkwzvLqxvxmoM
/omKTDzkxLUl6dtawO2VlxOBaithFHshZMiEjxs79th9qgxmicK29k077RSbABzrps3lQMbDS2iL
7Vx1KXmN08N0VPA8XPzeVH+tgWDNtZQBRRR26l78i2mJY9RKAyISbBj/4+9jANpZkZWiGJ83azdL
1CDVYi7skwIeKtR5LeBkC8yRIIFQbrmTiztDTdJcr2vvMT5t3MUVjA2rYhaVgoCvIviu63R3Xs11
4228fo4beqbBxjBcooSHEppRpe91Y07til7JaMWm8v8OjjuqqR6xp/a7ak0nEXQiRy2ayse7o0mU
J4mpW49b1YPdJYTQ5a2TK2nJ8qWAcHG6GGLlDgRxbcVIjRh4zcx3jE5U3w4m+pFdCgO15jMv+for
Ue5Pkd4smXJc43jVUoLPGA5TpT/SXNn9TG0tvhOUxS95dmMZOi093trmu1+TNjeE9pgwOG2vr7T1
HZxwRDyc8wAO+uqypGNwfvSaPg2LycP5il8cvAiRSS3Px4bE1W5icVQRGYGWrjt1zqzvD1pzfwsy
Q4V9pAJm2X33Oq8sZ66ZewKh69LS94mX12+ln3xIP0gfER+PHGQp+fxMOzv9dtNjCgvGLg2bkvxz
1ia9EVc5xNxIrZJV9Q1kk4CRM3hMDC4VpT3qr1E4n7qY/js4wwqZ3ASMlgjV33gBKFlrPe+R5V1P
vW6fVN2La6vqrigA8A1dwXZRtPOqYf4T26pXLJMRR68UVlAy4CV/MPtNYBLgVr+0WmP4v5jdidaZ
GI4xx3OjmQNrVX7rdu41Xu3dSWIzN0TV3yTLF97WnHs/aiCtsyyvav3FDQv89Msrb456phhMxVgG
pmzk+33IoHg/MdVSM0rET/MYi/jnik4TTJNa2kQdtMZGtN5FatvssH2S6218YG37OJeJspV3NFmy
AEODcThpaMnkYVpKrt2Amjo7gTjhXdfyIAZ8wBtmLeYt79WJHfkn8hmSi3hpfNBQKui6KIJWODAS
gP71Oo4CKsAGP5Oooeh57XRTDKCSPRncVub8ReuRjyQl6buBRexd7+hnw1c/sFSBqcsKL8nZuW4v
WCqgaNd3zhOe7B1AhwIn/m8R9KeRAIh5zlROAryo1UhmFSApMZw2iBfImZWv45XvJK7Xc/ycllJx
h0UjACveq3/Q+7NV6VMjK1eA6/KqJ6SJyEQe8UYYqDkhZVIhw5JntG8nN+BZSAUKb3iNCzp3c2Rj
0j8qjt6KILjKtnEED3+4qHfLLp6ujVAXXMxffHU9ZylYop8E7oVBfh3I4iL2uIXWOh2BqZqAp60V
ATUWVyLTaSNgdE7kU/BO2kWD126fsltQUoAz763M10tLh10hu8/LGDkHSP4VHriUikX1ewO+YPsw
jxJavmVQh3ICJGz0A3vUdr0e6zKrLUNv1lb42T7xW+7lPnvBdKk8cjqJRIm+jqs2STXQ4KzyB1Ep
fHgAcbunNI1Xg3SmiYebbOAdCFr2XUIhrCB6Te4kmc4KfoNdEe6DO5KsrOf3uqINjzq9WKsa2P/N
fWrXjGdfPzaYsbPeVAfBR0nAAGHRZHFOnm32jYQ20eVx1/qavWmwV/qYt3ktVwlTqeq7cYcjNCHx
pOUjo+oxE2pgsvsYdqsw7sK5OGRfvEVwXpySfs3jpC8Al904lsff1dOavN/uajz5OKO03gxf/RdB
EkuDqmLAiwxPvvT188LwAxmksh28dAl3krXhGJQQ8jQRUNm7vUA3mab0dQBkyrdt7bEBDZZ8x7Fr
IXBlSA+2g6+1hZOgruAplPNo9TZupQRy5c3JWBY9X5SQoz6IvHtGe25dBXIYPxTdXsplPOwqJDl9
IhTCTfb7zM+m2cC2zOXnpaHoanuDSmBOgwzPmyMUoXi3NJ+mo6IgCUEQuXvcTDQaDAtZ6PEvDv7Y
JV7kvfOiGHW7RWsy/1a6cPGtOUKjfNufAKzJ4HnKjKQ89UUIN1X1ely6VdxB0HyN4FQ+mXg/+//h
KF8ANavyFqWUE5iLolq7vPneJpqIkEw3PI0R4eon7Xa39G/V3BUSySkDqTxqc26iC1xFI0QeV6I/
ucpmaxz7TPvg6Wb74cI7swGks3+rWFVIf+yvg277q9WVj6taAGkOonUuBVlYHORLXgJsZaq7AWTD
dLY1yF+QXdV03jnSkclb3uCvAJD6w7rHz2jCuym6hyi9N34P/8KgQhj0URh2PT1NIXomueP1fL2d
0eCHlZrr1S4zk6KacSkSwGN8p9c22NGIraR2oeqKjNY+4QfG2SrpAaLGT5Sl6rJEM/RsAVb8ZmID
defRBEvlu3UnESFlxNlLzr0om0aeIds1V+KITzCzkEHO0O9GNcc9BR/aGYmlb5B0+6J3Mulmaz2j
VwLRVQrBG/ztSM0v4A9fvVfxzg+G8kIXDQACel983eib5CGOZVjVvKeDG9ausjy1eo0qq/UOHYCL
hePFyjmwByKEYMugBSpy7w2kRIBTtggPjUOAUm3DmTIB/tfb3Xn/rhM/rclLWfBiE91AW49tsH0z
KbFHGdVhxVxq3X6JJ1bUko4ZbvUXp3iHejs2JYsD8fK6wVx9f1YretZ3mo1AJWaakPvTSrCm0vY/
N/iDk+9+GaVuT+pcq9y8HovAwJ4+TZTHDjWXOppvqM8+n4rg2rRlZUtdpNA8tZs1pq0SajZG3yFI
RuTu/Rv88YGjTnBFaZIkicjG1afUyCp2ATc7pYBHz9j5Ftce2uQVgpGnhctlailxb08vtGqAbzQg
vTe3xqdWOULhgu3hUBaQivPw8HPMuRK1gPvpeX7ETnWNDQhUwLqO+aRfQ0O5BTE+tPO2hUVPR80K
YQYxhuWswET3Nm+81/64Q+/zN7peTa7zY5ouRB0+Qby03VY92IZwn1pgMoR3YI4WonDv6gKIGnKK
DLXW9BYFdvjyp0typPJueH0BXOsFqXR+JDPYM2Y3AyEIWtRgwbroS0Wz0RtiZ1DupoqNjLUUroso
z0qYN/Jf0/NsVtTqyO9tLlY0a+FZWSyfi6PLJCPn1mASMini0/3/KZ6BhSipCEPtsGfR2kogTE/C
jK6gWMeSLBtk+D5u0S1KXKU/RSKhu7MrWKga25eBgdmQYs0Enil/cZa2kgF2ldnACnek5L3ZblF0
R1HozM9228W/KgN2+FRN/dAWGbb6pfYUn+eG2Yz96AMVRcwJJXry/9OIm+KLlVqCI11qy2Yh8Syx
L6VrJ1DZfh5Qb0iL6qpGYkbjsrkFpjGNsbc90t7+Y4BPd9lWuHdoe6ll1By0PkVc2NL1PYEjB5HW
A1vht9CsTmqdJY68EhvrLKVBl5wLpC9a1dWTXYe8lNCcWZ3X4LUGeZ/AGsleCHhJGtvYUMa5KfvH
Sg65fLNM8FkcxIt4VNAzx5uCmgSDByX/KxwQi77SwwGQt38p7r5ux7BbRsqpxFfh7+6ywl3pnO9w
UW4v9CaM3nxQ9EJQmO82tcevWvkPzUFG2eXJ/OzL3n5o9zrns2bLlaNEg+ORnWiw+EgstUqy+Dqq
MmwxM24EBI9i6w/9k1vahUYDdGM8ULoFoN4IKqLbygMrOP+WJY7F1HQmPM20wnZJJBKMaIHRXYuE
lRxZnZuYVec5T5KrUs+tYZXqtJNvHf+gGBRB/lNxKr8TQuyh9VKZqecwqPjZnHYgXYKvHUbKyp9B
dpOW4kh5VUl8TC108DzWOYIMzcy/Gj9plC2SgJFkBJdMK/93OOL/89/2AiyY+lRjbZ1QvVNGbTAB
giiBOo1rUvuEwZGshE+/6jnARb17YZU5fOWWGWYuf+K2emKU3MAU6cmgo7tChvln3mTSfndiIKko
dgvXoaMOCw3S1PMf9goVgB+uzfEPlN5z7UvjZU57X1JLRdIxu+cuZes5kz2NooUi2dxFPz3jJ84J
t/CeVAmqSFdvZL78kn6wFE7dl1LdpnCH5oZ8W64ciwqW0HObxWW0BiRoUSz5aq7PnxNnVuP8iUbl
fMG6DQ1dUubAlB0aYtAKiEq3gHFCEHQHkiIZ3zapV/b5j/g2986hnwb8UvIOuhEqXcmCHgr/uJoN
oWTIRuIJ0Z6UbL8glD9fXj1bcgG7FvfsWiDzbpgsjPLmvi+R/MDsqI3AYTCWQaMmJ7VC3Z7OcVrG
qKKRdzD9VplNPzq5vxPkM0oFEc3liAV3RETU+gyaPbwpcEcxz5TwC+87yxlHv+Vg6oLhF6mOfXk4
qafSIfzfIeAlPAIXsiHCMsI61pLO3vy2ip5SdwqygbXcfTVu+QvBupZBESWFISPbkSd94OD6V3vz
/M2/n3QorKr82ecZsyBpWhlv4QlmU6xaO7rZ7ZQp+UQz/dCytMDUjuSmrw3tdDJUkc07z1plBNuF
eJD2uMEMlGgyfs0u7A39twdxAa66mUXvTsGMmq9LAoIrq4f6RIQCgkjMnZkMQOgxOhYvp7nFtXEf
jShRjjodTn90R3P2Wqdr4TxgU22EZyEKBI46izzswbdEV+yDYzsbKbPq2sDfOcDAGj8Wp+OkWuAD
Zlf9vYEzbjpgvYPbJl8j3NfMasGqj40hKycCw+HYVGY9rxSkhcpCEeD/fvZwL0UEb+sSh9nZWENS
Es/+SWREcM/oCmFCZUw2eYn6J274LNoJz761tc/w3pwz4xrz7r7NXRzrDgYewUya4Xk58M0ts2sB
BNh++XRIPCSmoEHL6JvCrzyCJ7fv/dyR9aeOQzT+s69vi13fyrxz/ozMU3h3RrL+VtEN0dOZ9wew
T/9L4r7tau9z9BYYKoaOa854biOY0ccQbFTAslg/LjeHn3dkRvXtdAlJ/OsdYrinWn+Pi8bSA9iq
DF0e99wfAQNWewlp0MjG9IXEs7MH9zZKpezIGY+8o5Qa6WJIvM09PrnUCAG0afNYxDCFYdsdh46R
OlO2dyDbCsFTqM8qJCNltC9iq57W3rH27eMKsBGO+gqVQmRn3vYj4dTVF+M/E4Mh3o3QQZXOYeA5
6t4E9ce+gbmCyEFTH6ABzVD9lOG1APcq30+d/Ipl4s+r4uiVolGU21CXwsLSmbTaYO3+aUYM7162
JiasI39hxWvm00nPtN/98vSHdKtORNwVJ0/Lr9WHNyvl2MbBhIAUmNe0hF464phEnmNPP4BNiwjz
PX+H+sXgJrfb++5IdxFODGfAbrkosrG+NHLdzB+Tgaxe6C2rvR15d0F9DwY/QFtmu7isNfUeQkRs
X5OP8a46K/sWKeHPqWYtnKIkxgYnhYgapYYGwGo/5ong5AWn0dRLQ1mucmLaaMkdhCRIamjK0zql
AsUCaXooaEVPdjUuoDhXBEBh1pT7G6UnGd9Yao5Xmikpx1XFRfq8yE/SqwxRJVyKPdhygksDqHle
dkLkexNFMQA4PTdnMpnPByLF6qoIMn2ppj+nxZuhB5L/piMOY1ZjOAk0WiVQygzFAKd8dC7SnE0n
z73ANsv+tBleLOgYgsRfZL3bfpDQreUfbUqd2ZNADvFoiQew326c2vLzKwJW2Mc+Z2SyjfQEPJx0
SZSne342acRl3stmNk8UsYiwkkE5sFzsswIqLSWg76w7Q1YTH/Bz6xVetCHuz0bVfsChf7bM6OTm
JMz3dU4rkn44iGIs+B9YWz3Yk4lIOty+ntOTcIr3bZ65+at1+aM4zfE73M6ov6lzeTspEgjBrguC
9GhjVd5ORz/d2nilPa6ce1nVQuNgHVHDK7JKVAt8tjbBrn2xruj56seQSvvrabpunfkRnXKN5n0S
SHukndWpeBWRmVSSeH/WsXFnPbKG5RLqVDXSuPJKFLLdCOMJ24POeMTAYjNW5OrkKY7tulWpKWg0
bUBbuVxeNGTmLWdH97qIbeWK7F0aTPxSJ2CBkRH9K0bE3Uq553BUDiWXq7grsItizNfUVGWZDg7l
KT7H1qS8OXaD8YMj+c1KWuzIWuDY3BZ882fV9MmeIEomdk9VXZ8deNxAVowsIPzx5hI7DukkU0Uu
1D4aB3ge3eAtD4ghqbB/Nq8pRlagb7H1m/CT6fWK9Cftar8vXMSif6eWjxv/CtgX9VFrQR+Ji4vy
akKs/U6tA0bWAhVXTOTaxoaHusxC1ehdecICdFzHJHMC+lSufniZNCV+QZ6tjkQZ2T5+vfzGkMii
n24wbBICtWdqQ2QNpDtqqmKB6i8ZuYBom9j3UcVYNZyp59CbwDmhrNly8wBMZ3SFRfH9k16mV+Rp
nWMGGoR4Lh/AArkT1nzORuoyzH8BQRxYkaDHKXoDO0aXfaVz3HAnq68+C/3xHoD5N5gbaP9qN+pB
ZNFucrkzDiIIVSLQxi22sa9mnNYDaWb5j4k8VnxiN2pwHvihZeicCShXb0NGXuTOv8xMTEIp6oIz
7ow4ZvhChXzxBrWrcjNuMxvlkY+ZCtahHMgvX5X+A/DLUwHq+UKqe3nPlDQxkSZ6Cw5O8mwpec3J
9LO8S4AT33Za2nwsXIgvc8UETm7RaGTRCLGX6Gu1lQM9Pw+HxqyL0eoADOThDjOUHwJD25sAPIQf
cq8y7rkyBdGxSnarIeUv7d9EmOHMBEXFU4DCHNvm6qx1Ne8qIx6Uk3lS2xcb1RgiIXTpAmfN0OAW
E4GdpcTkceTtZ1NkiLMfJvq4sfQsTqRXtTGjkQQ1GliE2JGb3Ea/pGooX7ZDZIXpu9Ki/lS1/Zsb
3fwr3jdiMojBD5KTpi6QwPaHJDoJnWkSFGEvu9jwpJt/Em+Ow3cv8R4gvWCgth5SmMxIKXC7p2Fw
2E9QmywXd+pUmXC+Eid+cNehCOs3a4+PADrpiLZuEQned27NBGqZtE4+F5F1NrgfTCMpTB1WS9au
N/FNg25cSAfMKAm0wM8LkgApJJs2PalcaUxmMAGoSmcVwJnHh4bVPp3GwUP5GIymXvArg4+NDLjR
DBOj7Gqd9WmbkYhkTfRkBKIKN2HHJzTfS1F+SYc3nciydXAVvv6S4FkBWJpgtciIkOwxOCwEnNJX
7Vw5ciJjDqZnytldHjSGN003DJnmj+I+Yxbn2fFIAi7xgNyLjO/yS/Bb2rYbp6KCmjNylu6chyRJ
9YTcORLTG4XC/Wa7Lah7fTTjyYuBT5GHLU4K0MTD9oKPK7xuebIulqNFKm1N84+jb9MJEXFF8qHr
lpOPErlZ8XIHKIAStPeujFZhkihynIYo6yU4VoIRLCv2uuNsts0OiLay6/IuX+A+KLTvbdMvVwrL
HlgmhA2KelzUQ/9QG23XFSF1qfWiBZNghVTLr0nZzKcikGdkfO7+d/Y1U/vP/RTOxHxyIOfVvBeC
nqzWk5fI/9cZpMgJXbX23xPqIT1O4q0G/TK4EvdRhlUrqoWeWcHMrLWPcSHIkwo/pKG8ID6g9K5F
ihUuk8nqEFMygm+zU/wB/S95YxM50VHZTz7TTsLnWefjo3YI88lmLKocjkmIxrWDUX0kRuPIDUd8
NzqGBbQHFRlkyY5XYSTLkTE1hnGeMZbVOoq2dodTPag8UP970WJCYNeqBcXY6pNQ5EJYniZsQbaB
7n5kWKZ0Z3E6E7e8+vIEGO+EFPPolTV95cN02fQ31yi1ZmOMFfycblWw3gOxA1IVW0fm1AKt9ync
/vSQ6RPMhhxdLRJp0O+vIHCYT6V/4e87qK50yUDy0IeqnGUKWYsbr9OzvL5Zme9ei8kUPmF7peXT
d040RxoyTxYkq0QzG8/AupdlXjwlvrGhDlZGKCGNEYjElICTCg/N1dt0Rg3J50gZreSY1/9k7M3W
YGID+aiGsjd2JQDA12Ay6aU7A0bIGMl3C/RLVrwzXXgDXd3ivCJVc2mpUM77curMXDs5pWgC3Ymx
5hZDO/fsJDr4iG0AOzROj3bVZ5Gux6BOuJbb3G3aE+Nz8qb9y8cA2DugZVSoMtCT6TEow1Kk90nl
dJ19v1YTrKFlBXC/Fu88aGceua9KU5kL57A/hpqoNeul87a9Y6VUziRuHR7uBJhvz0azDkS2D76l
6oqW5F56MLnM5mcqhRntnCylL+sYbcT3UZqav3sxxDLfThSUNo8QlussQ0tUrLNZpvQ+tQznh1ZU
5I+CAgnwH9HpZM9aJRY4yRykCWM1S0VpsD9I7ySMxN5s33IXhOrbp8jq1iw0vNvWhYsj+9PGAJBx
zqNvrSWExlpoavk0P3AT8+LC4YA2IYYb2hVloBMzXkqgLxx3w33K2YVYsSzzptQ+kT9/EJVR2Poj
ZmHJnnFhKoZZZ7IDLXVLNZGZ2YNSm6EFBg5T78/1aJlnskwfXZLXqQr52mhd3tW6A7jnsaBINmp5
e9qaVq3DCi1suqJYynmJwgushji+Rq27DVYA3fs1w0QcX/Hs6MinH7QIyWmMyx24Pt5AKHWOxgn3
7UIkTPh0+MBPdS1mWlJOMT7OL7EOrIqglM5YyaqZZROuKC+ztagcfyZovGRkpcQ3AGXKq5ZI22z6
N2ec/986oXQMm1a7sn3KN+WKABnA7e2kX8cHImjxaaIJfj3S12g4gSjALWrC2XADlfhQGfBG4u59
FDX6uycZaI2PoBKDMnq87XqPU4zrfZHgDX88uIYrKcRvPDPjbYIBR3BH+ykZfDlN6SNsICqkLGiI
BVPOkGoezvsgTzXGyKNfMC6I6X+uJatPIJVbF5E9Zxbf+1KHAB4qiDmEMmscqOIcVWszk1qODTUh
YKRjQBx5b1azA3ARfXNkHSpGCfPkYtzWtpreTImBy4S64QcKCdBQ3kZoydCx/HX7Ox14+VKNPRH1
y2hdEt7D+c2M8Vlvvs2GtA+8o5YFogDaD8D95dRq7N2DudEoJHrKaqkhLmgOLNX7vQ0+vEVFqH89
0LPaQr2NSk07XP219fdRHNKOyGDaAxAQ9ObmTN3Z3Ux8XuJvdSYvGr3t9e6osXQOHZ4HS4bMah40
gGrm7zSuGSLSSzM+ar3q+C4N2g5wgq9ewioQnoJhpEtl9+ELwpxbuXK0kQ1RW8ZtC13mNQD6aaZr
bA4RlOqm/lBHhDAXDPLDxQvO1ZsQ0SJXkXFMkI8wcmdsIIMdTLFvkJEYsKLvHuCp3bcEPg0W7ALw
vqe2pLQQbMXNXcUida6LXx49xefS77987Hp61Acq1OX/WDti0WuoqDP+4mOGfYsiC9NlijfVKsB2
Aw1YOYy1t6fGzRMwH7Gqn/Jal9U4w0ct8usjVjUF6RulyWnGgjTLncI9dBZNZDEZzP4J96lALVrl
PWk4mp1Qz7FJMVMzYPetFM9ZCTCxv+oU0aAiKQNNDvUv8a3jmC6MaIcrwfX6EnNG6n+W3kdeIIeT
A4gijw3MA36gbvDdPHqy46EGdJ7OVblI5Qa8ol8wA3Yo7eetmLwqZ7tyrnKkX1//fODiYLMgnwDP
CSYMYKByzx0prc17WUr4m8KGqt8mb4D6lWrLtZBlmgh8cXS9TZN8wqoMRAFEQbs/Bt8J0WABqwEu
VsZfD7VHaVRpwzzELa7wL0+IePqjP9XFhNxanz88EfyXB+SbyulfPVDmcc4QscPkiruPvuNn+t+S
znYSSjIZBDinDWoFQO/WxqjE9/TG3P/2RngCRpF/ywQdSxqTYNilV+S57W8vkRNiU9pBJORgjG2F
K3pmEGA/1P/IBz0VA8Lzcxlzn42GK/whD+wn7vUA95/NzbbULtBEDz5JH8RbtIDrCYI72wWAXjYN
/qR6LBP8n+MK79laYCcUQg4k65gdfpj5454VR706bx/yCoBsKzJfca6WbKpJQ0JOWY9T1Uv9GBe2
MnU22/JABDenHExt1gmRXuWq2NJx/DtU5t7XGZMVjESjHFyRQqMcy0eIdqA1gb99Retd6F5wXbet
qQZme3cc/8fYa+AVA7bBsU2rbcmI4Q1SDqjIGzQE7yRX9HeQiESvHLHUFLz6Sxki7VHz7BBS1MX2
VpFCCK1p2fOmmxmOecDcXH0ULkfC3hhL2fzulg2zD9jcvAg+NWfnin/bZpaO8Hln6vp0nH9LaUrL
Tf9LQ/CqdXOh5jWPY0thut8OdZUwDDnHadHj5qK9+pF/MrJP9i+ZVZEaa7CB+l15EdP7fkF4DHB0
Gf8lRGSmhktnKwDVBvfOXDogkGFL2yeGKxdlMxjvMkRh5vj5wY47P5CNx1lF7WV17zSsCMP3bmvq
0qnW5db/DN0RkBcLq7SLgQ9DsAFPWmal4jRzVt2PY8Z5cTZUxZ80xkoYSjz4lmlvkSl6t73L6cxz
Gg6hoJMO1PB578hBPVj5Y+ph1MNCpAIH8H0yFtIc7fuWvfB8Aa32dRNiazvvOwM0J45ZQkMmAU1/
xv76kr2oeJQi2kK3X1Xv+dL/fWZmJFOPF6Yt+7U/uticjwhe7sl9tuXrJVu8imX3ly8aRwETnEaI
DFA8ebpMj1mitrmV4RkUY89sVqKvAYtpdYEWgH6BGue+nImUIZX6hVfqCTUw/k6jZ4QMi0TAKFQe
L4j803adjYQJFQ7LqZcA0uxjwDz7DxBk41MiExiB5Nurwcd/CH56JtXBke59TkUkF6Uqh1yFXSai
pFJ4CZqFTZCg9eHmmVxu10Z13GdNMucIEJYeuRmNXDT+KagOaWsBnaLvxjvIlCRfUXNUFchYtb+b
Rv3NrZkuyHoKXnXSuwy63ehdq98kUYTyeBtHx+t1W20S8zFPmDk125uFGkM9uyhzVk+TaYxHrqa0
Ogv7+Bs1I2k+QVOq0d8cjCizSQcCqQ7gX9DjJT2xeY8UvUln65ikgWzCc712Nd1YPJdscb+YFum2
6Vqqtj0nPxrInuvERhgYY5eRsVako0tOPiQsI6Jsw/pX7HiVlrLmh2xqtMThBbsj3v+KLy2Fk+7e
HybjoSsii514s7b7LWLC5zqA1NmmQUfYHXBN5NaNsW4SDsURwGdgsT6NupgYT1DdyMR9yd2RlmDN
rxMgpQflAVvB7NSCN7cC9vVgPUsSZKkByVk3uAjuOBY7x6idQBldW5CSNmd0jfe3FLMJrojJF6uF
QH72iMPsecilmB66kA6jhUwuRzzOsVUFlbBLeFqKMWYmSr1i5/HmNGSSlcAJfbjll8a5Ys1hXFqA
P97Q/GDIWTU/VJFOPSIB7iQ3W8oXkCoEwxmTS9K/pH220qlfziqhZx/h7ekTjlsBvfa6lNI7ZeIR
ZVr5bPop4iKWGszwEqvFiTn8EEbGriQDhC0sCB5eAc04PwOJLosU7PMnWZlq0puCZVsQcGf12W43
cE2N/ZeJSdg4MA6lVxQdG6uRLesvVHaxGLtnNwDdgv4N0BULtDEzOkB3I2Q0wHiQkbpEyWhU3t6v
kKn/qg5LmocYxIHj2J7yAS+LAfSDRG5HFrUyWCa7aNya32DhN+/VmsPzxJKszu13XkRRj2nUmFzf
5lXOmbPmjxhKhY+0MF01tkxQ+CCfGvU9WGGglwpgzvViu27aExNuybWhXeVpVpvR2KEkLb1gG+Mk
eBJtggLiOoxpMDUtJDxgeGDExv0vjUWzIXcAL6c+g7i1iAw302xcVRQGFwaEXftE5gs9gAHGLOY/
X6kD1QmuW1sYkGg1J7/wCzPjdORSYJG7R+Zr8WHkXSIe4nO6VHkqP/pVOweMIik0GcAl4anJa8BK
Z3+G4uxSba4k5C2yNmqdzjaABMgdJcE+M2kynTOyFAR4mJUS/7k7ycIT1iniEizq5jAAgZml0Eyh
RMPGI3GDC1Iqmazdre0ltjUvKYrEdOR5qw8bHocehUlzfsLlictUTFQ/1OZpu3LZG1dRtkeGLkd8
BMFAKKqHtpDXH2t+vtxSr5mwo2cJ4CqTVqNjfV0YogsfwnjMLFlg2GEpEsg9YKy1wgg1b2LFUkTq
j83M/Hu1GvDgcjZXByv2pugzaEflX97TvTTn+LBB3uTtQ9VLRC7v/Bz/CKF7vYdzuCbWAP4PckiQ
yVvJg0s+RukyY0atvCcnpLXET/iraAG9w+ZLn+8nqgpsh06DoBHrmajiFSQOtfs1isSTtC3LlM2W
SwtPQW14tp5LwYA4Bwp5q4n6lg067LXl//zF5BzlCAs2EERIQReStCbVOj8T1heWxhK9u3jw/LQE
dLLN3+duKUb/ZbVO5h2nIMazuRLMFOetx3t+vTUhjKni15nuxTdoHvKVT8I46e2r3qDVOc0vRf+J
jfkI6gWnevGP4pmQi+uRDouiI9d72bhdJv/o7/n0sCTZ+JBGWkiokE7SAbX/BsoUM/NEl84Ipx0H
o7x/Wynezu+pgkxvaIl+lRbalkaMaPH9THN199JZeNWsJLl6pf4jhxw6Zl0lopa0isnnpsG6OxUd
LVZC/G+Zy4A2uuYf02b4W/3Ow0//wIWrS1eujC2nSYSZMDHHdd9U1cGa1PltXSe9nGXoCX6VAZBe
/bjJp6eE7d9fPMHTO6BqxaErjT0h4qz6M6CilNmWaQi90g2PgoiGVL5pfBs0xPgULk1VjXGIwD5K
oUiTOfmN39NY51PdAADUv7/gO93CUkldD/KNncEUycELWKtiFVk1qaI1ttICpKt5jJwIbStVNvSi
2+Hv/KjMJ5JG+LyldS9a5hX8GuhKMYX9lg4O9vdRHmdjIiwXaCufsFyDs9naQIwKLrGKRSSfBwos
CsrXDv9yG1q8kfVjNI+KAZ5r5c1+O8Si8vkjcI6iOaMikvWRYeJRNJo2JeMo/mkUZ0OeTHrnqka5
q+PAQgrWdiHGXHxs2EzpF5ApTlNyPdzRNHNGlHklSfqak1/Debn0ZPFkevpL6f44JmhOVdbLBJI/
+PQ1xlcuMqLr2XUsy04I2Qt27O0ZMHcsf2CB1rpxGvOS4Ly4E3ofdo0OslFZwWj0wOz5x7NnOQcI
S5uIr9E2As37qe8J7VxZc5hriVIhP7Z6yXADi+PrBAlVJ77rTJbP3Bvkq2pWj7S53o+jYP+4i0Cu
h+Ft3tkJHRTEYjCKBA5euXSvjDzBr9vr1xXoQm5N74KpCXVX49gLh/RafF9NwLTb/0W/Jkh1IESh
8an4Y8W2PV/rdujKBJ7E/awU422okIyVcCXWqCZ1H+GwkuGuh91qN3qcuRDwh4Y1BYRY3nJdOthW
/cFB9LNfEdAIMsMo+Ng943pLHaLQTpPpkjwaSXGiH65k5mwZFNaEwjSO35YjKjaogItqLjFvYLCo
PfDkpRXKdAWT8qCKOQeZNTOcpjVYYMTDAhvPILK/N/OEcTByB2RKQfRweqO8tTUiAMGXwog/VzXS
7F52RzQIPSPsGz2XFbRCoC7N8Yqsnx/0trM9iHvmUfdrj4XjLOhBz5rug9Q3Vod2LVZcVLKcsqyC
leA1g4h5z4vNZKTu51ulGjLPawLXO0UC753xoHDa08EYh0b8fgGeT81Tq23thiKD0vVMr2pQtsTb
yKZdsdyuxrIRJTrYGDpfnKOi7oB7EVsORofHAhSlDYEyI9yaoEuiyOdqaVBQBS2rzkdF/qKRbFqn
pGKvp4tNatcJn8l9BUIL2FiSJ2sQ7C+ourbq4kVqNNWmLrDht5qqZYy7lhFIrgtjKkPWPMV4tl6S
Tg5qfXY+COlN66b5TZt7FknosqO06Gp3kLLhpQ7yjMTHndq4nvtbY+QcCX2WAxZTamMKeNdM3Wb4
52kyzC9ZCT9iZTqzVu3ecc04B4Jnf4nnzGtiuxb6TuLtMKtjyWLD3eN9AHfB/D47ydK+ob9zCFfo
fALiXZcBNpNZ1mHlJyLvHua9lAOXRma2FpYfouoGMgiwDGAhQxbxRVNzyxgBD6rtb9uAmDcuEHdp
z+bLxLXh4xxvmyyaVvqP7VgCjOvd7O0bTDokI9l/e9egXYvb4qt5E5OTxDet/UYbjJNLe72MIaWT
7/U6Fp0zjBWvomOL91Zdfu6yMABY62bjyTBQr5lwbAn1RFjZpvDIXCKHL07DGAGcnNdJp6/rGtej
6WlK41bvYmW6jvzJGaumVvI5BSCArTR70KbMsBZ2mbWsM9tdLZDppCCSq/AUSOm4Z+5UR3LlqSAp
fTFQvhIfPvIdkpStE0K+CIfSJNi2dEobBbgLV7X/g24bTxZSuWA5JZW/M36S+V0pqVR3hNxcuQM8
hVxGzZ2dMYG5+6ZA6j1OmLB/B6SeRbIt28AGpDmp2jZMMIWT9Gf5YMtEdjT/11AEs/RyN4xcq9Ge
597NNMHV974aByu/ir11zefkeAES3pgW9Jonloe6Kh5k+OkNLaCVEgq/IzS4/OHfTJP/VuASKFD+
KnvF45lOkH2+XYUibhb1JnUukHb2h5q/cCufGcQKsxoPOppXdWOHi7Arc52RFmlevGJWNMexVx1W
lf5cKq/keexZ2GgkFSx85SxJ+ZNnPmXchuFXwLBVHHSWJPTQ8WYL1Hq4WWRJ8pTAxGbNhGFyL/lo
7E9P4VihxTDfUw1hxyhUMIh6N/rPvndrTRFFReqb1hmFiMYAvC4STJ/Mg0cS6aY0qhic0uDI7Gfw
Y7B/Nd1omkeFo+U/xXc9dRfXV0N/ELVTSymnkRUPpM1/1ZCj4iG+GJ9dLUdQCtlh2eT/qoL0YIe5
u0sbJHuVjH2Nhe2/GNEcgWuVsXfORbPzBeyn94bMm+9d2GVvLMLW8mTTZdJLGkj79HpmjbVlKRb3
8hm/P3ZHIYausj5AdIkBMjU5WxUhI+AMGR4P33cmiekSqV4Brmg7ZVMAqVJbJMm8VTpronMgOVcu
V1NYqdqKs2gStGmF9hJMstZSvyyN21RXkGngNL3TY1XeELoN2jRlXG64vN/qQMaLda2nZPGwoKvP
+8nkzoXA9I3alQoCcU+rn4a6CtYDTKBaEBgOy+eej/QIwaY+thgB7IbVP5y7Xu7grgjeqf9KwHe/
id/meZwZO3kPH48QIo3oIC1RU3ecvWEtuT+Ra4nqovoNnjZAWtT7jWIfRebqmNjbA0pCOXcYXr1a
uapeXIBksdsIia4j3j4effNZr79m7QMcpL9xVT+HWyqVmaCR+VA0ZzDVWDuOdJJv1DFpOpZYM/Ps
xHZ7FyemubkUXDe8QjfIbtLMRMTjcbBNnkBXopxmy0rAm03BdofqikhCcbiAjWe1OmE3w3F7ULtp
1oT8bmLQtewdIlNGhLfGzsrN7VbHGxAdljbAX5nkr7DMWb4ahHBYOf2s9vWvvKabvXRyYrFwz/Sv
GJ1cl6LbOtd+mOiFU52xVvlZiDsg5+9iARIxUZVkxsDh/ubO7L2rFqtOV3K3UlDxC64lwh0p9KrY
qGgzG1mLGaego/ulwnQvKZ0dUhpdzLrp40htAPZw8fM996RPQW5/sUZSn1UajwlQwC5+2UA3ceXm
gTZHXhSb4T/VarzrB5YO54HZMdW5EQuYXavZ2oGLMTnmSvdjmyW5BE61+QvGDu7f/Y/5ku3Z2aK3
koLUxPFPXctQRAWcRGMPpOwzuz9wFrPeGgvz8BsOcYDkkPUZYrGj+n15OxGrSzFYfUgwiJEqi68H
EJrHD2EV/Q2JvfeBo2+wnCdXfA1N0WgI60EEudLAVIBrHzUtTsNExpeIhh37qLvjrpN3UJJXZ6t9
uU3palE2xlBxoYwwzyXbtsWLoNW18MNeiXLP92v3PQgXhmUFozyJJReYontjoDhmpCLjnBWwaUl4
/4BuGSq94/juBWltu4N24W1+MLruLVBKqh9PLUTE6vSmWK2o/dbTkXWoHDTFs2K9cqbf01Le+fDs
K9svRaJ9bAkvCFEXKP7YVMFq8UlFs82hVAiP4NO4SivTmgn6GRdGIncfbCBrWk+ldUopaIoWUfMN
IB0buHLf/12IPhkOnHTz30vT55UEpeKaJo0pTYMdtTIX0U8ZOtr+wpPM1zU37VFbwn7PS9eTUBqN
53PkHKXha/1XObCZQOe7MdAkravIf1WsK9Mg7QDpfbOCcnlRqhyH9sonTxVhAz6TjoWHduiLUVf6
nqw9Xmqp1gvPi7wKaejPhnvUN4WAQ24j4ax7UQBqI35Xhi0BbPmndP77DZo7Hv+FeT41cdABF+FL
PTqay9Q6F8sQAkBWkQP6f3vkXiNXrA1jE03vbsHn1a06KHhTvbQbjFhjlgV7GKMbblT3lBRjZzYb
Yj98lyzJaVAspcM1hGLy8ubSTzrPRQxcLTTMVKN2DuNQeCf5A5Lj1TaDFIoYi3RMB+RkT7xTn7SZ
60ismBbgXwpzKrpV4WlrmZyYc8DX0gVE0D7L0LYNby2kWTBIklFqEjqZDb1bf1AL0YQfTcvlmGsq
6psT67Pl2lGgCfYSfj+gRMMDti3OrairaKX3SH3r6wXoKba8u70p24dN1KtZLQqLZnQsHmlTu4a7
ROUwHnUG0Ld0ZiwzxgUJJ/rZqH9YNIQhrtat4RSuKfc0kkixbFW4Bn63BBQQSpWY50INRL5MBEeT
QOU46pm0p4OPK7akO5bGlaHLXD4S1usmoy9/U5yVcIqystETIjsQ4MRkmNXFqPXHpR8WJX7zDXun
jAxugzZDMkfFHKXUgpNPTejsgmAUHQiaT00BZ71pM2JLUiVxcqNfOg6BKyS8aBc9nrJOI+tKYOZw
yVSE6+UKwjMjeHVIh1ywrzMFG5yWSENivG3PhYuQCa3ml5JeXwvFSfRXe1lhFr4vBMuOIBjCN/o/
tHQvSsEtDdMW2avlm0ZQ7meCeLM4IBqhH3SyXynNnN88v7MULato4kDTTnhTvYuEsVDw2+BNxg5j
JkkTQQV2XbVrzLcVec5u44cUOr15Z549UJj/ri0+qQf6yTZgyAXr5jwFk0XKROz0BpztBuwOt4PK
5z0QZ2Nw5dDZ4M97MU0SN3vU2MlIWAKkOqCmYfuROpoM0UExBRkDF3gsLYm+uhKfNFjXIQdTke9z
J50fraSn/jfVbMxBHXWZ4UYfDEwrQWFPkyfBzRQj5xmiSzc5dZngKCOjiVRzH+P3jzaY4TbrI9HT
10SSA7v4JuTb9DbVgBV3v4Fnj5mFXiPqGNC4PVKwCByBCLFUiMmNoL4/OKKFTL6lws+YjWj01Jws
YPMVpFrEFkFZ21fnOZYAekhgWhK8oDpZrsMJzzaCrbVQoVvuNJUjMytZAH/k7SPpkwKsGhCy2v6p
AVxDAuLTeS146uFApvCWTq6xMgKWqgPPnUnvDQe09IfiOL9mrNduJ4HJ3exIs2l1Deej27ReP7XP
BCD7kIZ3uTBOdhO+fF5pKCyVnuy0sKiTnhV7+Nlip/YTS1rzRvxIaKMm6FirzCiZCdciyj2DKHSI
p7TImGcPav5JR4zCx8cyaCYfpCw7LiS8ECUmnoXZHjO4J5ibtIML09T/azBBJMLt4y6XZp+MH57q
f+XKxQBQYf0vwuqiKMOA7lpvGsf+MKKJq/9l1elqqw6EWESCmHytBDtL+Gs48/8/lu5bTA3Xd3db
hGlDv6qxW5Z0Yz4scrsXC3MTQ1MEcDl4Uw35Dt30e9w8sX9n8KRrLLqCpdCWmyezE3FIjluehg2T
7SSlSxl/sHMcLmXMWWIlrFG+0UZPiTwyUSMZCEC7u3d9gOsvKOy+W2sdvwZ013hdl3we3zdL3fqL
QBjYD/tTa7mY35E1lmEhrSRq+khVkHyW5ow0k65yEh0tHT0YugIC7WnGodPzEu5soSr0lqnuOYTG
umeq7acORRa2B1j8rSjGpY3m/h1tEQ7AMLcnZBk2Z599o03hn5C+BjoG5XKLjpqFg2IC0oAjdXHE
vcOJZe0sIY4qXzefx0J3YS1TAUnUkPfvqTitgxRPqteWw3v+DghXi+3t1w/WX9PmuB3xHNjAT1jQ
boovYIkC6/wddW/x3aUgK6IkKtv20YohgRQNYwXJ0rqKwEShgfMnWCFEd15yogRuXbOL7sMfQJeD
pWcJfbhfNe3bi4YfPGg9dBbI8MLNPYuQhdpLNGrSmPB863TLEe4sG9sRIF4dsTG6r//pET+FTgRC
6pcMJTYgbc38YAR5amHYWjSbxdIvw1Zjd6eQuj2ZiVo+PoBVKLwKqG4NDp2vygY/jd/Mh3afQMfg
oGOOa9YrbRmiixE9CpYb1lU981qUX57Fy634s50uxFu02gAQTw40hZuib+yk1yF0Ry2LSl1jaCSZ
FthpeUxnhL8p24p2peoyElYq70ZFjNDhpnBNPhpETcpyF4pUSJPrji3HkR+XbcMKH8qWsT/pxkuY
y37iprpv6ZfKqkaWVjRNBzgvkA/DVspW/zd6iI2Xe/XkAJf2kmBe3oAybspRnQfmhEn2Z7J2+jzD
cCvGMSgzixafJNOxouVMwFpvBI+Q3NhhcXskEDygNmqLHm9bP7i1nPX+NKPP+cAcVeLQP3AT/Iwy
j9q4KUeqYHdfzi4Xqkb2ijhRJj1pVGe8q30PJOaL6m4kfR7w9ulzwrMKZgKM1PWn9K/r5ATh60EJ
muHBwR0rdVgmU9DWwHMw+WY+muZu/Zou5eJBJjmG8tv2ReQzrdkEPDYOZkyrTadeDSASGWayhWQs
83p/EVBUIw7SYPqZUE0jILRkmfNFcvAmK+hfpkeZLtiR7VR5eIaM/8A3AoMWT9uyWYlD1WoFKkHJ
y6jAx/RCW3AbCQy9osg9nVVzbIBp3id0gIqxwTmeZ31nAYwse0Eoygilh1iUZRBFIrtC1EAnHXpn
GjE7jG1OetzS7bLzuQ8geG0+OBhFIxmB3X7fdz9pd+C76echeLgkHb7cDiRCy115FDsyXqSc5CeF
BYlhKdWOrTi7o5zbRo5Iu2rbqbFWjaT2z0VG74qhI8pM5lpYlfsj95g5LGqcpCPLZj8ITyFYbkO4
f2djM6/Q4dBl5ynwXe/EcqrB8UleLVHVUpYtG4sN7PTjMeifWWx2ZuoClvPd7gLtFnF2WzJgynvc
a0cry8dbPjckjINrE3h1fI/s/IKlhfwXsAJfuoO0ZxPquaAaU+UD/u/WLM9i8eYVFhEEaCwRxJUs
F0wcKJdUZCyvXn/EWEyDXgHP78RHGIYwh3IG2ptM/15BWFtRVxPA/+McXUGwajWoiclUgl0fw2p/
7I78cSKgzC1Mqca1hCRAGOg7dms7D5N3jg7OKVyPwtwmy/zpTRhVyfWdZiixfymR2Qz+3GSUbNYp
gv65SVvZxBRVYWAAoujDQT7stZRnl+XILJlureamtwp2pgFChgWykFI/sTO0O19U2CPmM3OIJhvA
rzT0kuk3soDdE1nN7kkHpvuSmpBu2ybtFhj5k8bnjZlu8GAQaSvUrO7Rra9pjwcA9AnjqmkEvcuD
lhFREmM8qotqK64U9fz4y24p2ejCVler7KjRJlmiCFTT9V6okUEIcNBpgb87C36SPGh6ZnRYG6M2
qV8NASnUkRfh5QBWwL/0Tg/GRtFHgTJ32AxO9KKGoTQ86J5uoQozSBWJgzRoeicGs+SpYxJ3PwtY
Jp9If8TEVYHOkc+INfpn8nkgw31SBxo6zvGfyDvMjlXvppwSzmOH78RFcy3FkzlDgZHEYxhRK8kd
mnqDDBGvcfO15jPNyyEHj3lbsZBoTHRrJRRsaRoQfdlJN+fZ3BP7SJ5EgAgInhqU8CSq0UzzccqR
Tv70EeoX6BGrsFG6p73eHUZSo9lLPhS2SpmI8sulXcCipS/wio2jveEt9uiRIrmXFOnq+LEEZA9G
rz2s2dXDpB30tGWQyihanqBsVrNyxuUPuEe7kJAI0Dtdwz6jjhqfLueseIiTqZHfuXeue2y1NhKu
OHUfhZhrBqkZ/DbMl1dR+LobonHbHIBce3g/tGs5kH3JK8AzlbA7/R8MBLIqihS2TVyWqQmftLBS
l60/GWzSah1IdBvkCGVif+gBRfbwtamVobk98rC6k4HE7iKJ162poDKTy4WOV895CF+H0WQdLNQE
l5X/Siyl8c7JDI0fDQhUw8E2AYdcrs7jovVsszSym6+v5FMtRdvrKUve/pBKW2VshwN5y/ch8MKA
ZxX+Ae9MQW9TSDrOXxGxc8Q5CZJUkBj5goy29+TUSjxFjh53/JojEmprZUlCfG+GDFo9oqoaBbV8
fvToSb755EufqNrLJCQpufI+exSeZ9jdwtyg8ms8GcrrV8pxlhcSLuHRfjgJ6WA8zEK1Y/tuL2TW
jbtlIsHx8FORf+FcHuaoumjKaG8HUJpLQG/u2HkF24+PEbqiUxXk/PKYF8sxN4OrVX3QmJgv8B80
2G0BpJfd3MLR7ooaA9c2bopTKbIRaeoN5fAyOOoLYt+U0OOMmtcuhcVct55vRCh6jbo1rhSuMa8Q
FCyW2TXesCbCk2P4tl/nfNH7hhCpK2wtx9oyll5lGtZfpJBqYtMzNJNFeFWtg3cdrwJ4AZvtqWP3
blcSlyJnWgsk6WKcq83uDUx8lRwDCW4kAeByi+g6hvfXa+nHercwbmQLQmEhp7jmAXbsFvTshcIR
8/78kkkSikfxlBkKJzggLtkfIaxU/pI+V3yXi1Pl197zv5YgZjWMM+lRNt/rz3ybDjysjsNZwDVh
L1umGpcBUA9nRzBgfaAPG0BjDPLfg/ZL4UDIe6wRxJbGokA3P5kOVYarUGojay6B+BLIxU8seqMx
4gVXqcPUEs/tU70fHaQ1EfIHYPe1F/fMlFsQtcBx4i3iuDb9nCsREvPGMg2ud03ap65o7gsWh1zN
s9cz1TYjqCTdJCMRYgXm2n5UGEn7+J+xIbM8kS6z2aBVQ+l2lhM3d2hWO7aZHknPQGZkQva/c8kT
EnwmtAUDEt13kqhBkEiFLIOZjp8xBFBtkd+7Ix2Tatf6OdzZWtlcIBK5hVDwKmV0EGNvMH5aoHPo
pkDlyPotum1CNAz57IV99TruEJhteBXHAGMM2CyOyT3SE5lx3rL6OQQlW6GMwcQREvZxo3xYQnDS
RcKtaTjVd/lLvlaPrf7M/lRJL+I5aF7lKT+DphPvECDA1yc67BKfH/TxiR+wKAehKPGaEWdfsApb
N49BDd3jXoIR5gKNIn3pJkIhcDC9nTaf5MY6wxx+I3heCN7uR2zcrvRx6/afzkwO3qTwYjXsKTZ/
BTMxwz8CfN4fsCv92QWpRyTpyoN/FlNBcCMjZ9gM2fT1oFbuVcU5FFKdgNkdEcsMLc5U8ABp9jrW
qibcK1ISV038LEqX1EtbemM2YHXAGUpdhglINxd7Ay+L6ZhKnyykwHfT31jfC1kIKrcgdpxvsHDb
txV0d9/w6S1ReJS14Pryaabqh2O2ZlVUwHgsf1hLVi++qq5eEr7eV72ZWwT4i5zDMj4KmrpqxY6Z
gje6jTM4qEkLGwFzS9+zcGupa902TOjKjVcW+JsJaMsgalp58lHjwFg/qzEh2u+twUZrHOvcelgk
JCo46M35jauuUEWeBbrZ4anlKM1UwcYfq5WvagRtgFc4okkzGayGsnpwXi9vx1x5yPZeuYSA5Vcq
DX2YblxOpkhNeGtIJRNmVD74a7UdwmOaNHJismCXKeLywXB3XXmWBEFM75h4yd+SC9JpL2uDwEYz
xom+3FZpoIUtd4/OoAvip3yNV52Gx3F8h/hPcmteXC94rvnpK2e6eGjESKmc1vCYhsM9+Y9KhoV0
U54Ht57Rei+vHjnYTJdLkG2Utoj8O+CltcFldPWv53ywh97bfRDqFqpGycaHADN7HP/QcgcKbAEp
VVRXRMDVyrCW0H5rWiw70itLGs6PEs7wBitrAKVS1RS99XLbJg/JvAAe/sq45GZ+ZSNdeYQ9FmAF
8EWbRDA+5kDR0XsxBYGzhJtiie6vKu1vpbjs7NTVxOKLYYiujIKQJy9bLIjr8pAU6RDat7+ky2EC
YAb7QhPWQSeWdyM6kRZWm8BMVImICrDyWJuOwpnRV2t6720IrhbCr/qSz52RyZULXoEofNZEumJ2
DUCCYq5VPy86kQp+OTuKIWnQIHMZrUn005TZrA/klB7WIuLcmYeCYJB673z651+vmouq+MX2kfR9
bh50nXGScGRcPv4GcFXgzwbWZElI2pkMCLE24vqd13D5ZxP0LzGZqU7+LsUeMv/HIe2Zd0uzCN6M
6D/cqmxpY4pbh1B2RhksPxsiVM+Jx3CxK+vpkdMTg7wrJ/zhig1JGTQUn9T6el9MnFIIRVa6T34R
3wpUcioVvi1MAqWU7svHmRzaBOlMx7oTv96RWesaPj43E3xn+m7ttZzKWr8s73LdqbPeZApcZ+3r
nl2/7yIIRidY3jhD/3EpVWVh3lAhCLbNrZBd2sMuBIifYr2KZtcAk5g6PQcp5y2QoGv1bl5eqpMt
LwfcU+5bE+D4bRh/d1P6cgZWkrYalhPntwHDY5ycWJgZEd78Ofr8/ubKDRZzQPbJdbVLLXJjudEO
sHAETuEy4yYXEwUTXutlPGAr77tSqD7X6LpD0+b/SVlqnqqe7bKMZsW77QUbo7hg0BuH+4V8QCMP
2Yd05g5mvTWVU3z0xo26hGfcCyU9jr7ukwkD31tRBHrDsJExrsgBiHyUEvQyL++gqabxV56RLeQ3
wwky9cRIU6j1a0kv/8iAzWaZZZOiyhJY/P1r05AfRuNWEA1dyl6pvc1sJMXofbpBsvauXEi0/fEa
0OI4q31eNdq7seCY6qQb140xORh/tdUG27g0r1aGmFOok1bL20mWq9YwZ5wcsNUi6hJj5WnnLWw9
qd+mrTQFN7AWDQZHgnEDsol1sqNeJ7JsICln2F22aZ1oSvUVCaH0lxz8R2E5yCigG1hRsvvFSxjY
iKRaWezgrW6Ma9Q4mpqpIT3UX3MZEwB/9x1lwy4S5eo+bsOrghR/HUFttTcOZdkxrE7hOHBaM2Gl
FoIej1a9/WkaJUwHHk7aF6tdbxJgxS9Sp2SoP37ETuVVxLG2dRKEyIkysSeMBdb4udbnwltl1nR4
oZ43DdlFWd2AvrreypTGd7L6A5q78MUXsdPd5LJzlXij994CF6lstVj+Ma+NUMYYRRowANFl6cFo
PfH6WGY0cH+wiSBc5KIB8ZzqXvrGKF0GI4xWYylDUnRbf0V8KdxmXrF1F6x+QwHAIU/6uy6dQyzh
sgj4qCJbx57UOMeODFiZVeTee2nC4ftYp00rSGJg38r7C/UntzfuivoWXd6vbaBAINJ0Zfb5bzDz
Nls5SmPVOqcHLCgWX1gZxb3OpnhNAURYDaS4p6CM+rXZLHZtAIDs0nMdIMMETAih3/gyy16TEddS
ZBoJg7DGn//NdACJypdcMU6KXODAkH+nJiisNNf9jKao/uHwUpDesWLIqxmvNGr6lh3qN6RU7t9D
RS7yn08mmDg30C4Bthzds8OSKdnaTx0dIU2V7xHM0N+XmbqiLGey2J5FGdDz49cNDkajIO0PNDTk
adTnflutv1V6x/59K0hoTtV34xCDOqT4Zrr0Jv+5w1bxFviB0M44dcI58xTkE6DnAfU+3fCydEAp
mnH2eop7apzO9jIuCiwW3Llfygcb/Ltv4YeB8u2Ga5mUmrrg3xDefbBDM6yv7o74KjtoC1hOU2zE
ty0mWWOKSbBFF7/EyN69ikUG0QBmsYH4eDqNCiVqmlhBG/VZQFf0mUnyLmebbD2zOVf9ABMkKMzo
/Ch6m3S9SAbRDJC1gUWV8UZOHIq+VI2BeuKrS3XAoxHiD2kOR3kWEKXciwvorl1D2JX58zjmjrej
TLexI2XvwHJqzsmZMugYc0vcPHEpiC1TMzwdHyuDB564geY9NAq4yeYzcqdgyPjK3dHOq4nCBitz
KJ+FvN450SrqCn+iJ4xbxUGNsSFJF9K2qMcgexiNuQImTmKBqUy+hGoBR6R/5yai23ONF/fEmAgB
x8dyiWRUD4bSxxe3gLrU1lzl8GPifT10ZseXb/8APS061MATQMFFX8Rcw9DwpUjS0GwstiFASxNq
ss271eDf1tnJbZ7AFGB0OpaDzNl/xOPtRZbDdSjk3yAiKx4bmDMA2Tr4Tv8MwNgArTZHso2GCj0f
E55ag7/hZprGvDg934+MIswY/FYAn1AixKCGm/syPCTRAkwHdBLMsYj8KPojwwzHwOjIpFp+KHhN
b6UvIiBXLVmxRPrn4tWpxX1YgWXLBVQkx5PqrP03EBsFGXCfKU/DVFY0GhGPyNqvUOnjIsXqBG9P
IjtjYPT4Pd1ZziKePbvUsgo9K9vgSm0WTgBGQ3L/z4xP3gKxn1UinnJvZ40MjlnbhxTBZlWq30Gi
oTurkcXYSUw0jpsi2hYLxjNpCVq5s9KmBPNF+HtnCsemWznygMbI4R5KhfDcAWSA3MfWxghHq8kJ
QBC/VLxyciO8NcMYz+V/2DCqAxJSwMGJi03HFZCrCxDpeMbjfkd0U6DrVTvXJJao3UKm2nhv6Gfc
5ueoc+gLmF1fobUa9FuPxBpsGtJe2KfG2JCPmXMAJMS/u/Kr/TBykNtQsTly2rq4+yPyc2BOGOft
OaWAqb6MYMIsWgoJnDKpFzbo+TI+Kd8FqXgFULnUsOvGHHG7qofE1e9FdpJ+H+ASSYJXHwfOmXML
t+XFaSPvt2MsffEaiksXR8JH+7tRpcmD/bOzxLNnPhCd6SRu+h5OYBkLVlgJwoeZ6oqxe0Ye7eAh
AcA8NqmahVxN1wD9jQUZhWWwxpWxoYLUoYrCRbKHYeL5296fj3ChrSFNcQpknGlxbTnpEItNzMtM
t/CfrGm/70Gx9HMJvCj5WMMjyWo7gfpViRbFHockIzWImisUR9e4GC2xfS7MPgKqniNGrr8DP+Af
t0EEyZYYrR5TZHueDJ8aNikVfBHRgtwPqxiIlcMGJyFYNfGN3IVeekN1dVTq9q/duV2MNCAd/3bw
rkN6LtwX5GCtay+3bEJnTq9RqsHQWLRcXJMm9w87iOYU/+zurB2CrK2wYcfalEXwOBAA7TQBD2WO
Q4O+2UaFqlOWw3kK5/hUr59XWnay2TsNE5sW6KwGRf6o6+DK/CxE56gff24LnxBZtrxDr5gPngku
qXf4Fu/+aTcN+FLshH91O7rF2XceOrsrk7FGbLG5K++CZKFLxru+2Gkw5MizVTXlbMwO2p5j3iNK
/KojRYEteCjJSDv/Pvjcrn/Kamj4OPQLJHYxLj6BujLjQF3uYEvARoadaO5DRzbRL7Ogw8YJno9P
MGPlJNCA0I+drVtwsAimSaZPws6lVNnoWWuQl+/jBsMmc5K9o0/gdsANnSjnoiWnak21hTiEd1ab
1ra0BdC86MA0uQ/SBQFpi5K3CC0eod6U1jczPLtYH9nOV+kZ+iveLSy1t7APTCTPp3TAkxe5uWSq
Fr5RWx/TFgSl6SYbwQsJEU5+bWSc7ZXydxljTQPl/IclVyEHH0L1hV2UJptIP7tK02OVyWA5SmMy
csF+rI5gdq/AxsMHwMH8lwFF1lRB5OapV8F8Lqk0p/tJ4lJ+iPcJzZ7E7GnLDrqj3yzQr82JawPV
BYuVzpegp+Z5JcrHRXd+ukCe6YxKPy9vBbzeM4FrIDJipsrJWxw2upDORg6lajn+CSYimr2Jt+wa
GwO1X0m+z/1mndcI8wehB2BCsnV1FJg2Q31vl9XGtpdxuT+vXobO0RxuDMSDdJyFoQtz1meurhZj
4t7SdprlV3ekBd2ikrcI1jJ4ZBrDae/OyzK0z0OzQUbmY6wbQcPobsCwxZCAvqtQ6/ikjWhHq+Cx
A+4lDAErSzTvYyi0NpNviMZ4mFMLgGmHh7Z5ycwaphlc8tCpDwF4qDv9ujcouHdueIwHVM8o6Z2B
YmQ5aFgrDsprNyJEAXw8SXkBCppSKXHq1vNEVKokq83BFtmU7pxO/9Zq93jJtcMRShV3a0/T1p+q
UlgSrMxnpKEX5wc6ad/QVL9WAu1N9iJp0o/RnP+wX6VB2bFRy7fwqVLO1mOkHAVXb+WKShgBjxgB
73FLuXhrPUWOUz60UGHkxVmchgY3AzcPTGRrlL++pqoHfZ11LdShYIev7yL5FWpnxz6BH09GeHOO
yKXE15crLL9BWDRjMc4VfiTZ1rx7d3H6w6krlz8yCJ8pBaWPgjYWa/lGRZ7Ozj+ktRtEQisHrVgh
JASrIGwnU382smHoNsvl+LoXmw7xAlCd+GBqBGXAdxBgLsK1l32SQ5s7wcxCTKCyDp/xe3GsaxXp
23YlJ2Gjy/aLCsBj6i+aK6YGyku02vjHwmJ3vae2lwKLIliP4l6lMXt7zrwOlJb/ouW/f914Izvv
FlOgb5NprdesvY8yV/73+Ntv+eRwsHJWM4G6bcb0oVw9l81UwYHcfYrtaTCLZEjyxwDHLvh1ha1c
uWHo96K/n/YM4gDKKZ89od4q2rtIB21cYk5PVH5O3Jfqnki/GeMQO81VJrReqd22b+levLiDyfQh
ZKNnEwBzGrMkzectMHXsHlEvmBNEgqTrrSSj9ay+70Xsu6vGqeHFPJjpz7nSBWaDeIiwxfa1/hm5
fweeW7Mpm9yXtIBIQvNBxY8hvyyiDnXG63bJUmn9baP5zRxqAbhyNXo+APAE2qttuj9dQma/DdMt
z6SLWY37sG5RL1fnNeHgAgLygcxHDkjscgVYDpeG7rBvHQhZRVX7CLInbTJSmPoHa09xDa68eV1F
shLBvYHwS5g0g1SPUo4qAW4iBtrqCVlU5gGHDho7ur5qBr//409zUi75HQK1oNSpwY86sTcgw8FZ
22wZxRG19XAQ4tXYZnMOfyhH69zrd7hSJUOducdsMuidJxVfJj/hNMYOp4Kl6219uK1QF70hzaMo
jpoGDX4vojK3eNFDW6ZosgDpfJZClWH+GNCfNObLKK+AqjBRec98r7sZIJXK2EiZGK7VHot56FvZ
9XDi7EguU4GAGgnbUI5djI5P3r1OPhz5qmI+me62cDAjOmbX2NDRyB0vdkNJ+8Cue5s1JwGQh+z+
ZfGcZ4b0H3p8AdSyR+7FynYxwRz+1plLxFcadkgsue+6jjn+dHG4PRbvJF4gbVwoq2hqyQejrQ7K
eBA/fkfNCTWL6p5t5exxv1CyucXuV5GPKNA0h/Mqed684QAZTfKUYMrWwtjEcgTHya0S3hEbtFDR
voCvdKGEDWfmIXKSzAcVYjqTJAzzoyoaqshCmQ2Etivv6/Gp3RJMPGdBraZsvx3fyXEz4xdnQdTy
utojuKdgaC/FOWBFkf4JegpRMN81dTTT7D5AUk1Oc72Q3tB2vO6SZVzouRj5SN6TGB/n6WcORaiE
HT00hZCeebrdYnY5j9klot+o2K0+OtUbMSxEnJSh4tyNk3OmWlPoS5NU1M/QdKKOmQ/1J4qSDIF+
aXt6YkrLcOep0VWnQOPYEKIYs1IfsJbrTrajbFGxyXF5+Bz6ZcmlxauMgORX8PlVNdahdZUoV3xd
hi9rlQxHRiWddjSZGJMr/CBhHgVLyJ7r+l5EdLYkszZtzOZD88/G+Ir9htLobmr/RKMquQVY2Rqa
yaSG7/UDKhzzQ6Ws2IGrNAyZa4fkntVhxNwXYVm3Awq7hSN+RbhegBsJ19THjTuIi1hJuiKEUyB6
D4Z80au9krzP99X4+AyXyvhENL6jg94h23eM0PbbbNIZAAfRlMQuyZX/bRJ+IuxeUyMVN6+psfpi
rH/OJzZFKn0TRop9cndC+EJ04FJUcYXaOnEdgmPhztaYrD/bt3QxSpH0E5D1r2W6GaDXBUpj2cFm
raC/IxX50FgodDJPDnLwpdwCVGP/61BW7apR+jK3gWQFqbqQoUCFl0kS4iWemsAmt0VUS9l9sBWF
qCbXk4fGVrDIMpViKFFUPKh/TOcuLWBJ6QVSYpSqpGbq8SENNtOfPfKq1xDDcG/LaJnI3RFC0b0r
ZTDkQK4KxQ7HDEraX2uW1byZZCu6f0p5uDIXWMwbegujBdm/VvWzyvmwwRRunu11x/HW1JziVGD9
N4cDwQMHsCZcBbpNtKQYiWxcbMO4B1ExbvIj8eVOiikwAHi7UDI2KfGgEgzBF+4nFvjjgWlx/dCv
Am/aRBPg8KgI1q+UDv/FgAZPBzv6FgYIuy4dyqTiOGINh+TjQxTq69kyjTC7nlROc6qXwQaKaFqM
7tshKGqK883j4r88VIVJrKiX7K7dHN/cxvwPBdTJqqefytfpuGV3cbPGJlfZTvte7o2K7XMEoGXY
W/pHI8/268iHFFubo/Kmou0udMd5gKk6a6FCeqjFafJJTunRx/oGIklZvUQ2elCK7ENp3Zh0MJRQ
vx1f0iwj4p6jUz186LRx6UxGUocDzSCG7GO6Lu+o2sUwv4VbvsCgtg7BiLN92BseluSOAMdeqBAA
nR3zZh6Fn0BQ4BSox1x98eIvJQMItn2n8ZgSWQ9/fTMn6Khu/l4G76M4h50WRvzz/Y6QBVHi8PKz
QmaBycJvLjtqCbNmKZx/8iCgJMLaoR//R9Dd9OTBhwUZYwQ0TZIqpOz0pyVRQtWePgGao9Gke6tR
X3o1hNXoMVTg8ztYOjNZ1pIte7DVjgN4hhCYyxtLsYLUj3h6vZR/7upo5kwDnTiG2BRMv3TabfuE
glv3fVhdVrf11T37GW+q48idFPDjkXgkTnxx1wJMZ+EX+DaytlBXBvUpiHLHMLxVGexk2cRZxE+a
0JPQe/JfIyxqdWomaxRh7mOEHspCc3a9hmCw2HhLAosJpCZGoOAIkVzKqKsaHwr9WrEjP0phxmVc
gGR5P6TOToBMc++f47SRaOtcCN3pDpoonAJ2tnvU0bBOLCFgOVZ+ftbAaWNRKsnWi96CUda783Gg
6KOiw+lxJbvHejEOj4nihHzLmWa383zZPt7/kZ32P8/KuAv3sl2Q8eXLt/ZOGK0lyG/q4NwtiCi/
t8pcKK/fvTq+ZQTlDaiMcSFXXkNpENbNc5BHXvYwjEuQ8QS5//S8Dt0KEOzsfi4SL3qi4mKW70ti
J/yAUMOqgGGxGYMHIBkmBqrjnyazNFSc/glU7lQU2XgzgTOyLM5TzycRBBSYZ0b8eZ45qPedKzv0
lfoMvsPogYHbxTcGeHeYCCAiuqiqkdWpFDz9RMz4KooO06CaofPh8h1VIynE2Nj1IvIleY/A9Loa
5c0LiOL7yXwy/2fSCAG0FZc6rvldvvg1d5UvOanqrhjCmrKEMY0uQxtJCbN8blh+rwCSHZ+xBMOl
OjDdPhaRLhNYv6Lo0rWGhZ+vO3ZYM+8hgdl+oVxrHC3GydJKcdDHiDpfPH0sqhDV1RSD6EL1VSnc
7Mt0suk5IJbCiWw+eBKKR9iHl1cnvm+J4aOPa5IB9k6sMxqvdnUG6XJKZQLO+L6x7t4XorY64+aQ
HCJq3OALX2nky1UECI5RIbwSx/6ch/59TcFjSdt0ULEzKhzoxIsusoNcd40UsNRo5zREJZLgLRdd
i53piQwYgd7dqeaALAnqlI2wdyHtVdMJkU2SzZhw6752WsDrN/2FIK7azlFQuzx53CUv8MXL4Vjm
gl1GH/nkZVknhoABXIB0aHDs0Hk/JJcVDVfgxg7auq9zLdA68NR6TFQMEQdtmdN4BrmRzHpLDgRQ
2qpN0f36mRkHwQKnuoSU2jNd0UA5OQKDVQWvqeMvYU7b+4CYSxU+Iw6EdRJwxW0WHNBoWe5o82Um
qwp8643QM2mgkJqQgoPq1t1xQAV4zfpOMk2bQDRBTMKi+uvfiz6bRXfIRDbHGJa7a6IxfB+0fzvV
e8Ax4xS+hXBjGjV4HBL66NwLG6RkzhqxgdxlR43mXDKnW+aA5KYGr975DyT1Qkar/a8hdJgfqpFB
PYnEkFmQYRUVm8N5acJ0sMCUVg+Cy1KO4CM4ZQ7IFVtOacAm38goN0NeRpvV8IaM6PRQCJNpYcGo
NGCKmpD+vGhpULt+ubp5nWDTTImo9gaMAnj4Na9nev/s6tXpx6K5fPg9Wu0Zzj0EuAUXQ+YFSi+t
bOhHnvAQrw2mtB2rznayYM44Dt3rDGKpSGn1LvzfgkixY2o6qTNc9WAqxmMbYIa+opJBN155rvO1
+lN6axUW6H3MOpACzvBFcgf72xdPGSMHTZaTdHblBGi2a10Mz9f/dvyXieuQ2dTbwDQLelaL2kPC
3mvwI8anV4K39/H9+tccBJwagVTn6KqHxykJ5OK4E39FTu1ZGrBDm2e79TuAQ0wbCCKruJ+OJ7TX
+sTjKOFSt1+YwRcSS1/68JiK0YSQYwNj089cQvNiIsBPYYpfeP42DX5l9hYB1IPSQSCnIuwvbJmM
wTfVWOrNGYlGRyHL1CLCqNsjuxxD8w0Q8z0gUGEC3hve4YP1z+wAfCpqVBNapJ0SczJjv88xLha1
/fBn+Et+cfNt0Uey8Q5ndlzo5gu+u+CbQZYhjhEdxIdjw6DkqKoc05VBZ/1UO2V6shTG5SJb7B+A
tyOsN0zCJZs/Hn+0mgijRqT7wIVCM5v/5/1I6ZoGMX15Dk/q6IfA3iR6yKvMkeY4s6IOQEE8BAlm
ZKEU68HRapXf7gBvXNQQQMOyxA7lKhzKGDggOpO1FHDVmIT4HFPXWUi0RGjTjtYhIMJuZQIVIf7y
4ysJvTE9P7J10nhuXHcmhmJsA4RCj8dIRozeEEdaP4CXm7XM0NnXqMQ+Ow580CMRT+onuyLkuSN0
bVqcJEhtx04yNKf2ddVkAhjQ6IPL42hSVn2CPOzG0/xvkBobkiQTSJvkrudL4CfWXgDa6KZAe3cj
Iuo3cD1+/42H41kzqfUU0b1h7xn9dAMyXpjkedCq6vTIqJsKF7IV7Ptb2Uar8JpuoVnqnW0dwA30
x5pWbweGhmDC88e2saYLMvY8M2npv9ZzIJxaVq8lV9lhhzD2uEIFONCDcfpemX839sVb+speX/qe
G3HsOrtL5U4UdJBPAV3LiH9A5+e3X9P8PrngvoYV+qED2IJlwMY9zcubybHHUu5hDUexyBpJetWe
nLXO6sHFx90/KOPYHRss2DhVe2cjbQVy/5Q9D1q7boTJO8hwGihIr3L3vjRWO6RnqyLkSYHzI5cC
LVblCp/lAHiUIZyoQLClnw6W5f+HSI4PMMU+suE4b9QnZ1hkm9eSHM5RuZtwz3hekuz15hsYsc3Y
6IGwS4eEHN74mT7JrRa1Vm9ac89LxBF5zFCkD/cusijTK3KH0OFaTqP50wFQDeGFDG5pswveNtiy
VKw38XJ7LYLhEGHkKSW1Nr4AHOTYsr6xxQ3TSnnCtx3UhDsA63jFNoI8pIu9Xufzp7zlSQPGQozN
5dqbYb3oQrBL6ouubAUqwaeHBRmLMNPCppGzOTs0FmYkr1iDVuaIxMNSi5Imk2IL1VGTsJX7T0Qu
iNwwI/34GW1Zn66Q3Pw7bpulIYl2eEMsFEaW2lJskxzLH9fuy1gv8X7KnRnJ2QXoLAkGh5N40j8l
XGYYoPHPqrse2BHeV9cAuMUadhO7kk+UFchzRXaeez+/uY3oAUJT9qZsPnv6IdfK1GZNT/VYExxd
5vGsqmyfkWj01lhsivMIlt3yDCy5fUsliLjLo0Lr1EyXBe0VIiz7cNAfL0p5cqBUHKJp3nMCChkr
9xDqd47JSUrZV/pPWbW97jBMP7Q4VuhJLjgi68UwGlRPgzHqWSVB8oo3CHamEFB7Q/BlWpQjdjrE
ZnT2U8y0euRESejK7OOsS59hD+VqUTuKyh/zIMbfqADJgSQf8Kk31c7piHiiu+MTcq83idKtqAz+
QGrx8K3zS97udKBwOnTRIDJEJok9cVasF4daHbJ4idf5GjGpTGaOvROtEvqXzjIzLGDKh1m8WFPI
+PP739X/TFYX25Dfr+0HEtN6asZEeqO42x0VTQOCGnKpzS8bGYt0olT/snD2THKsalnTHWjqhal3
+1DuvO2Da/BT8+Noo/+I13XYFiOsN5/dQ4JWjwfP61RXRDT0nyzq3qs7rV89VuWHZhxUsjDv0VfO
WU9OO7usPuGknaQdLD05jPY2BJrb4MM4sKzxbYFNSpgGjq3zv7qxcG+MraCK6eW4j+gaWWrVr//g
r1GGGYdjGJHsrbEb2ORH5O3U91YH+Q1JyS/CnL3brHEX737zZvLc8OABcC9b9KyS/KBpdFdkZVec
ZqfINRxzDzqx+HVz1qDeKso/eioZJ6npuIdadpEtIpQLNUqjbuwTBwuCMKgbkOKEBl0dj4gDa3Ft
VvlXZ/8xeNL6rLcYgrn6mgH9XSt6LjxWGFHYy9/V8OymssFD/YRhH9xaZTE7AVyoPFJ9xcP5FeT3
nPGTPKS0EfYyLUNzFGP4+ZPQtY9A903Uf1Ngw/DtO3IrHghE0yUWnLM7BoZC1Dlt4IFI9TWKl2HO
h4i0yZ5nixC4jSDKhXZ8xD8wth2BnT7vGBzasLZzBNjHVfGFW5C5tmYy9FKvUXV+Ldv5DAsyeHQT
gkZLv1W06SlNCv/vVbLtP2hN0GIGiWtLlLQLouYzpEdRq6tro/SYePlbf7VVajL/rQuUFHTt8xDx
4SZrIEqE+tqFn37gM4rKtv33r4d8sdhD4yE5aUiQ4nm6yZ6fGA0GPMZ8w+CKN7/IuTCtbi9BsIVD
8SUfE9CeV5T9c+4ijoBXTvjyagMO8VXPSUUwX9b3jIfgwJEzRsTbKnuglHlHYCWRADu6zbfpDLPr
JVEy9tlOLwone3Z31MY6xpl5FNzpetOG3QfTeXU8FwPNST92h2vKVYwSMIGulejTAdAYvwA6zGkh
fyUXxvur/ADWLzyVBCgi1qCC3QTaHort0ymUoU8RqwhT73/YVYaguPM7JIvDzk95fWl1PQ5ezP3m
eaejUgoYz/Vckz9eFozXYix+mJIgsyb42RyMdKum9Q5IuOYD3s+x0Lr/rxTmDn78jjW9CMCIGrTx
9C/1LP9IE6nqXEwe9VIXClCLmsyZDgaR5zAIpCHZqR4TA5C8YIBXYjVAQFXsynRS7VC8cyH17YnI
XwW+d7kOEyn/YGUCfsJGh4V61ztRnwMtTcM+IRw+QHBDq2Hq6xeHPLRUCpx1ldOB6+Nc6xZ2ypo9
KP8gxGBYxpQq6FrSEj6Xp6vd0dFmxeRoXNwO2RqyKaCoQT8EnkqFf51RVRGGDVd4SrQMBV1yF8gL
VWSaPLf2AJ54j6pLyXkmB75HD/G4OXxVc661C6kTtiUlYqo85dGZWfTPPR08RAyuReMGslb/7MaH
DBjvNCdE4rHUrGne7y/u9JlLzT0qKnH2xdA4qQ1W1XFffBHZwC3YzbQKJvPiLoY2Mk/YmXfofbV1
jjfwvtYDNjjABNfgZncsMuInA0ichG7RaLju6apiYsIbROd9N8HG23WlYIzLtxZ6Jtlx+minLDfc
zHmkidy5PkfoEtMKXhjylB2G4VbBsaU7wddlSU454CAHBYR3tsPZ6HrrJvl9XRaKdm8o3uzj8pZa
6TWlKq9y+rD0TkwoquzabFGiFkX3NLyXkdDh+v9iCqqrxVdHLegqgVlFCk1hgRSbzBZ9nd3cS99S
1osONNWpBPA0Gm3rZa6BVHoKT0j3uDsdV5wTW/TtqjrnKlQ3mD39VoxsHXnFttybIbNRe0V7KG62
6xNAviRKagDhG/vH7vD0ZXzeudeDRY6pyb9TgvCJTGRnpvsUfzQWeEtZrRsI0y1OdyCUXlnyyS3B
LmnSDER1jDwDiGDpYvLNba1dXclCm3om2jHzHQTFS88AnnREaEqy94tUFBiAq3OnHJ5ycA2sZrDr
Pzvlaz3MI70YYof1rKTO30tKsqBmx2AhZt1xn3nSF8AhxKc95o9Wu1SMdmh13SyYEOwzep8pzPLE
ckH4tz6qB08J1ORUIVwYA49hyTNeheDM/jaL8kXauRYRreSy/UZhN31xe3H6ynojGxNKODkpCt9T
FimDSTjLtHp/LGFQq/BhvV4G8U2FdgfYU/ZqVJQa0f51b6DvEiUamRtD+mM0DaehGosjQNtvQop0
gADdk0yYQHGP1qiHQB2wi/BvIwLr0+3svmpHPnvM59f/B+JX2pjpvztx+0/OVLiu+8eO9oEHQ4/4
dE/P9HvK+/tjivzhdn7QUeOADWmSyv7S5EsxchoWedqlL5z9o9lpmQwa8s7uFFfWCYzGOrBgIGje
OMJXbsJSDYIYzRBbtJdnrwC3Y86Bn1Bz7LSYPz2pcGr/JpXafvjVgxPKHzP9X/Rd/ilP4dGBPH5a
kj76f3b/MjfoaBJqohOixJkRvsjFmf9TQR4wAMqZJ6yYH+wI5Wx86JrcTE2xvclVen8/NWODB2MS
ZXD2xiK0FAbvhuHYMkDDJIH/D4zIARaooSlhfPQM1h8Jiu45OUtmu5i/U0iXEENIJ+88jTDKbVa3
pwH86lzCAErRlu1NTjJgzfBxyLck1MEWUmitRJEOG0liEQ26K68T7s4yyoNkiFAFQV47FwGqFzdH
lcpSXQPhP4T1Z0/8bsZrPjIy8cDGEP/NH5hMaDH9qXH5o3zGI1tKZ75a74DU1LSWVTIJ3N0ULXwj
qHzD/kA0oMiWqy8DD81FkD7gvjH6G6xJhOyAN8BgHrQEvRguUc3LWpiaw1NGNI+vMK9E7gjPkMC5
DSuSB1gqrv0pfyX6uzN0UCr0/7quoAn43kAjQjSqdkwtvnV1sgwtnk0UHWdKCRikn15PWEtY7Zx4
OvW2K7XDN17yj6jdMi1rcavnEgMCT1LhP34ZiSk/fJbtLtrxOb9C1l9FWTb3PM1wfLssmdSpzexQ
S6al+xOSrGJ3fGUhoxRWyTZyw/CwaEk1tFU9KeGALSt/N40b5BjrgIykRl5mhDR3qWPJjyeRTIXD
CPnxgLAd25QNScEPLRYwA3uLu1Uu+ouBnYt5dlxu2xii6y7K6wKJSVFDe04r6DTvJ+keZJyNdA2V
Z5AcIOgw7+yIgDjQguAF0mCjN4+/HJFrrGZrpet4MAudapPkgMANUkvbI19vqFxDXnnKmnpUKBkg
komQf5iaX6sxR/njBBFqIIhCS996cbUjAiV/dMF0dwkcqRno8d1kUbVoe86k6zoNX5WV79sGpEzS
aGjGGJBWHksyDDRqxX/Hvp49ZlgQvS5e4zAGUoQiPU2iWVCbn7zZC17vk3O62mg6A2yJAa9WgbqP
KUs1e228KuQLdrrf84h0v0qur4RArcQQqufyhbII/UG6UarHglj0CJHlJmL7DjqPCoeHQFgqq7YK
Rlmz0XnNSc+Syp+KA3ZPPMXBzp0xzSXuF6/EgAazvVpiASqw/eZQoVJ5aBkQtJRjvsMBuAmrDOMK
p2kOfEYgHvjcoQbw8Wj5JdXUnB9yIKqQLOe7awdy48fT5/0sZ2QGnpe1fkNXbJdteaciBn1ZrhPv
tF4jI18HVTknoe4t2e0Umw0vB5L+4MW0wjU+L4a/qR6LneVx0+OwjInw7v29dcMQjMSLWAgT6SMM
1l9VnzchpNrsTwgHUgo+rVEf7H4Hw1fLoeapvMhYN9QA8ssBLxXPv1aaSRv5RMONe8TqNJv3LaXQ
mAr2fDjSLJw+Sy9BkmsDVBT/c027gRU4+knl/cUh3d5jOYBumGsbtFKXXNN8Z7aD8CT4UpEPyXoc
ZyJMTYPOYUsauS0saVy/Tw4ooE+aib71npKd7UiOnBN2k494zo61fPMJ8pPLsAoQei68Vqrl9v05
q+JA3mKPRmsYh/dH5m7rJR7WgZxtRHkvoGccyeXbm/ZEFdX1+An/xzDp1h167lClyt+TNqgk9CwC
3k/UMFz5fi7apCJlHXa4AdR3NKE+i29IragTri2FkAjEYqwTvYvBQZ6WKqKk3zBeGoSQmWtNcjlM
juaH90sJt71sN/eunOVul+uT8tz5cMzvYP6RN0hKDDIXmwB2wxqWjxqilqkRy2pc2SaFw043mUlB
02LLVT5tdHE2YoeBU3Gnc70LDGghKfShfpJNNPdwBu+60ZagzpaiwnXLqPoAp34bJhI3NFeBKhdN
mrAFeIOVyhY3OmykVSPRWn3EEdnstLbrqo4oofKl484mL5iZVsiff0fM/R4ihy+7nKYK/mBsolnj
fuuMrBqKQlrrqqb5O/wbrofz4HkIVpKfVQlMsGcygDJBhAGe14w+UgAFOocSW8cNgzyC78qNq5+k
fyNQCnOHI+TXgzkS2yaBjsOjSurlsaK2eAguZ03dzThWXgCA4QpODHddNNjoW16h1gzmnZSSr4XU
oQSUkWnnYzCFQva+fTXzelX/ywmgKfzqgPr+Dw7D35daITmhcon6s7Pw/sguRiVQLaQC+YTX6MaU
EFrMKNC5JPS7XeVS28GRLV73lPRlVAZAX+MQOt1UWrS+krAnNhxzHe4KYvamK970h8JZ2y7lRzqq
urhiMO5gL4lMwIjg7SpoS8omQTHkKfG2rkZNtNJOeG4ftdHwPIOWBNpMespN3REGbzoM7WSIrEZA
fXv9LJ+bS3H1M91apPSp4NfSbrh/62XXiEtDiXQtEqOyefKfXzYlkayRArsN0uwcv+8SN6d4KueX
2yoqNzwiRENE2d5N/upamsrNNXqeK5NAj2W+QoitGAjtoxeSsjrOTPzyak1627yTUPqeiCdjCafi
LAP8H6Ht2piIAmPO6uXgFvFurg0pdW+mi2N7wWhwZoo5iFyXnd4AvS99eDifT3ZjnDGF3DOCeCN7
GD7wjx5RxxT3jmJuG3SxniQx6sS3SJXgiAlyPK4T0BNmun1ZbTXAVJLtSD35LQ2AxvbA25yVGRdX
PIbONXhaIIKzDaN5ASJ3Jf+9o8AxC0loyWK30L3q0/TfGGf3xi4SA+4QpHucZZZfKuypLx7rzqk8
VKC6wF08ILyMFhdZOubnys4OdFzghhjcbViwLTDO+8qizj53pLvfBY/wn5t6rCWqXV7WEiVzLWOF
HfszK+/HjFD3mfuabuzNmvSzJnTCPOxvSXr05gB1oJHNrQ8SOUhTd/qo6Trcap1p0dh7is2jyVoU
kcmTZwB+rLhOZLS0pQIXCSvzJ8tXZZ1w6ZnEyxOM4mRHir7OeUouKUGXhQ2ib4c9oqme4LIAp3Y1
EF2LnwzP8Y6yW16jq72FJwmyRCM6T24yTpJqt8UK+49zbBLOaX0gTDXz4mqEmi6FGo/T90sDjRrf
ElMXSuQClayOTXK/gymF979u8BMH9E86ADCQMyTHMgE7kd53FVJBa/Nf6OrItXG+rAelHkafvY2i
GfZtRTOEE1P9udJ0bdSvJNxS+opdoRGpY4PltO/uKzNrgEv4s+H4Uyc/AB8eY6yOOzV3p7ANuz/T
FgDeQJ1Toe1spM7vc6JwsuwZXOa3O2fqPB43L4sRU+C4311DEIoi+KS6KfylA66pA42VYFlgx6qU
jDaN+J/jjjauUREn1nRypjiL2pj9myIlSthXiMTdagTu4cD1aryzoABMWtAUk8CMaCMvgsU9wcTB
7qOS7yfI/zvC72cFdeLt+m05Efb4BSUq/Gzakj4IXUn95Md3KD7S8leLoJA98CA4kH6FZeKY2RSd
JgkTzGcmDwZ5V8iuym70YrzME+sBOcHBqqnBc58jwGFgp/qhqsYnQHrN8lq0OZ/Ejhll6PNPI7UI
fNJrP1tMIjlt2AG0HiYJlRE4uMUVWGrkx/miB2264xQUmYUKfzE0tulboN3h12MJMxxpvQHY8f3i
f7GyKM5qGQuqIGdsRgNdlPkJHBBep88zE9mcvihm4QQrG8w0Yr/sFpfEHVef/0AHz8OpMGsiJA6F
JaZDVW4pbk5t5ArWYlJNCQSjzdUh14IIvO4IerV/FEdzCn37uy7tmTWqtEloyvh4JfNXSeGNnued
LCZicgEzjQZQJWy/Ckl6Y6Dw14CXCJ4gNlZaXACvV+qfPelQh4+85auDZoJBfW4SXr5L14U1JVDE
MBLS+GSpVnJcDjcJwJMWcoHFp8gJdv3e/j96rYWMsCeqUDu5k28BhF07qc8td/84WRKIFyu8bNle
6IDVVzrXT35v2DiKHFGyQG22AkNndaS9SQ2cP2aR8hJbJTnfbdwRMHdy83B/hMqJBw7whGaS2KIH
+noEZ06z76u9AqwuAqdxjWGO3VXB6+VaKINNYo8/4oB7UdJi7/zsq0OZ4X5ItZJZqVDch0wPpYx9
GNNDEN9VB6MK9rg60cqJO3fafho6L1V6AAF+HbXINv1lZpDdoEz6VJ3UEesV7bf2hASSsk/sX0yT
kCRCKnu8HEh/jVaqZyHB4xAg0JLzl6Yio7PdePDR/2T0CpNGs90VORPlkKQ1CDbFXk+vLm7rMvC5
vI+c/l0Q4Kj2ksabbz8wK0eF53tDL5qXUIrqkwlssur7b+hfM4aCUL5bgBlxGVwthCuyw0oDbYc2
BaVdia9l9v4/obr/6Q+JZc1AdpxQMlFnJ0WPL3Az/kT8Mcdj7E5u2AHpjGhRWs7dr14TGQtzDuje
tLT2XKN5M/YU8GHURNgYDUjIPnZZ42abLoNHdADlmB9R0GGnGgqGdGzsyXQXE4zbb1QpRddGiiut
Fp2i4qat5AVibHENuqSte64zH2HpIgzAopJ81yb+d3YmBtDrzGjsrbhIpxxATh4a+eZc7glVTlxx
6xmDnP1JHAzkExqUS3bSLm+bl2/XwmnVhX1lNh87HMYyb+Ngrwy1DmMUMonWJIJKuZnzI//DKiPz
q+xbUqQInuZA0la63JKn+u+WAK0WZC9E6HnFc1mpbLLAx93vHwyE1+S/h0X08xRZUQ70N6Z7+HXz
lLVM5sM53sG8NYVXC4vVfRx771D1Vy/ks0nOeDXRJBH1Vvd4qzzzlxKqOgMsxGcGBM1SobL65+5k
ULpDHDe96HJuOO1vfobhGPfdmm3i9McPVz1CtTq/a1uuTCWpAo+tss9p7lJlzj4GUgtB42uAPqFP
yzbf8JbEhNKZV+JPDOKI7kPYyftHpbhsAKX/jTFt938Io4CZxsjO/mkkltTUOog+i6xMeFR6IbVS
BMqxlN6+CDDVwYQKbKqHcBTURPBtQnfe1JIKAbgbEKRuBpH5eLRO7pJovK0jDPDoQb5txJ2lx1t9
wmaGMDGJlZRcOommNlh+an61OeG+qjOHFd7vjlaj3avl2VYfdXxh3d2/WNqSL68Hp1iNJGEFeNS3
JDFRFDj93WbZFjaWHP3/PYE/t+Xb/YITkWUXKSKQzdQKev1zcBMhYKfGAGWDZQn9Zu3kY9HDwZtK
j6WdqgvqCwPMCGgfiJddkqkCpLYvWsGvporK4fxQS+myvgMZFm39kUxBqf27yotC8eO3DW2i7Xjc
Heka8hw61oNZQkVcvsZEDSzTubWX7y8SBkeqZEKus8GqIz5ik4EGnPblX/i0D9FCyGBFWAFccrlS
E+Fzk/pjUFyDPPvNF2WvQzXPomFtzoZdhWMFLmQAOg/z4x2NqFLDu468yh+mwf708vkuIwUowIq9
XNfN0vj0lKOOjkCZnB7cHrwnGIav7U91o9f+qBjUFhC1Ef9y3ICpiqtjI73M+iHzbxlf0Z8QP7XE
iM34TppBc9ww3p5dBtW2Nuea23ZH9GPf307eNIzwOHwTbXwgSIhA8u6BNtNt6rq2eGODqSg/ugZC
nzPzP84otTm06z8TMzN0pNnvhIAhAYnjhyFsFhoGi5j64zFRR7fBQ0KCIGLzgYJIEz2De1W8FQg3
EXdW1IyBGsR/nfytj57uLSOgQFIkHwwHoqsC4Aq6cR3xpBsaZOCAvCe0D2Vv6J2xPeq+hBsVghcb
EkkdAI+6JeL/5kT6cC7ckSDD66n0/jJXZbxWZWIBERLgu6oWSuUF3/QevGq+++U6Fw7KD+P+TC5r
gn3I5w51ZrpWFLriD0HKSdaTqgSqIjEEFr3cpYmlAcqtc6D0G3fJfPbRz45rp4wNTsIarSU8wCQY
wl1ZoWa0pB02919RtRvYGrPM5r8/jxX7E/BMrbgvF5tci1/1DSoMbu7YsVivL63HD0e7zBqtR2cO
OC2xCVn7CMKbpJ7Pve+C05FGBf286xF6VjP9ocZb0zUXgPgcBJ6AjPd8WZnFm6ijwvAYqQpDL19K
zsWxFX+TBLTuGiZA49NlEr8Qv/SRvtSIo4jg91ORge91b96cw1zhBw9+d+qhGpb/g6OutH3X1v1g
0QB/FowrtR5Y2ib42RpnCmPAidyzWrm469aIDmxPawbUBisoOLq7chqUnsxM+l9luThHqEU9i/gS
/a06sLk45Fh6DKHP6bI6l1k205gK1ug+UYYXsK2ACHu6flaFzF/hJvM3VW/GtfitA1RfGgwhplSa
gWGpLI+U2q4UHLrGRIZeaK+WDHD4LOVmre2r/C2oqSE4Od7Sg9I3gMl6OVVx39paJRDJo0JWYqPh
i/z55+Kgwi4DDdAMXFhEkAFABTR70nNylv41oTZqYJLfkYVP5LDHUzg/mETNfKy9Tu/dR3RSekiq
12rkxP/4sgoVKYM7z1reEThCN2/dG6VnsBgDMl2F7u0/tnWfM0BqGibchABH/K4dvfRmEnhHPsT4
jfdX91hpnjX7/cvW30F+Mz+BbmbbaPl08qEwV5Gstou8INQ2IfsLg1BB2y3ogvI+liZyjZ/OpbxG
eL6ouPB3QPJX7PUBEvk59g349QhrsRY/PX5fYdBUJsMcDooMLdi9ivtLbqYXVUP2zcu2F4HdWAC2
uDoksaZy3/tYYFzOhTmG+GY83ZFbR//NhU5zSiH1PiV7LVVdsC1JYrJ405bZs8/lkdTv1eUzePyc
4ph02+J77gwXy70drgVoYKiXSpwEJZ9WiCC0Kz27uAwlIwMoIX5pl7oDovVyk2Wz+RvupVddQhfB
nOEjmrc5j6Zi9Td8YALgqXeKgHdOwsqtFesR6XPmQaWPZyETGtdyfszjqb1uoskwodbrFV14TY3V
3MtmBkrqUkHMZnSy4Zme/N4Opdl4aWdcCvvHQWVA3MUyvE4Z/nZin670kzYl2sNbY4mZ+NepP+BJ
le9MAziRgVVFHqlCL5N/dVGe/vEAKruOC1fEUCrQV9mMXpkj9NmhCAgdCZZHonn79oO9bt+Kv+cY
X6qoyO1kjAiN+dbRBQ9yenftZMctZ+LEi++xQPColCUko3IF/Z15lPiAzxSWzmid9/j1GiCuultV
aDPj1roctgeVhaiCAkMPHYD1cfQVw18XI1YQ+vzotvvj4EDV07O2rHCXNwYaPMqaLeHCOjE7YNLv
hh2ygyMP+uXGYIsnlAPODWss7X5/ZvWuMAAcB4V7YOzPgWZkVRjlm+dUfWzGqXaJhBsODJFmGR5u
hNva7zYxhY8vRP/9BP6NxIg2RGNtVLp2dF87pMB+lZq7pinaSTMgIKYmr0spje5RMKA95v7ij76c
38zvLf3mehNMgI0ruoZaM0uqvDzjGAD+ytDc4fbnu6IpV8FsByiRdq4GByBEVu9svgS4lBq26vOy
h8q7PpaD3NhydN5LkZDHcAENjwAZpUEhFfyGl5nOGB/8PFpkw7Rvqc/2592JJX/sAYH/+8DLDOTG
X6i9SpijFo4gDa8IqeTali4fngdEe8Dpllvpmhan6PDHppGpF/JSGR3vXhwW8U6/myolFhh7QVWf
cdGq2o3QzhKasFFFxG0vQzBEr+9mQxNkT6vsTOwAdzLt6DHh+0ha15YEAwmcd0kFzc2Dm7TROEkV
18MwSIbl4YBG9CAkHl7uYIETplVwbk2g/hGQKv6hfk/AMSUTaSo203TJji+iBkrtlQH2xQ2kqtEt
kK+J74NyTGr+PT/qCPZ9cWI+tV1r6J0Qz5Kz+h4+uHgTGQV40E5fJrX+709sy7/KD82A/5sKVd9u
NlU/m9iWgEemTDa4Xv0Zwj3qzVkVVDaaNljljqUtjvY9a8c6T7ivmZEGdGa8i0loMcftxkGnuP1R
PfwXp8vbieL67+eSqqTRjpBKWHiz0yQzaom0MkXy7Ogsizbc/Ysm882YRPSGW5orV8aNklFMRdfp
GTkoIh0TBmcDBvnN1uIxpd3cvxepn1wYDE093mhyOIhg6ldeZZFlTilr+5bZ6TaRtjXZrDnICFJu
O9bNK7+JUXqOGUjuXnX9/eRz1ShZ9siI23pz35ShwS71+dGQNLo7DROz8qvd2epWIN3TfHP/e2vE
8+G96/PNx3mS0MbUvBvxpiQ3610GBG/ENYybeBiq9iYQzV7g3nHLTzzrZGSUh2fjGEfAKMgLkOcW
awSYE677KNDrABeWtTxEpY+rAE8X3xDHQHK8TiQ4jb9fEGPKbObqjNOPpdy2yoK22MJNHcrTYk0t
dktOLLoXoKymToIf2cwHDmmRhwEYhsicAHlROMCIMinVepDvLxmVRJTVLSh3o5DPxhHE7H4RBj1h
Cg/9+sx2kk8bhJLJmrGe5Qns3G/2hYNbRm6sgR1Y3FZkDpYKqSnBG2DK48VMmlzU5qFxk7KaFPlK
JNAtKadIFZ0aJPiaBIpgj9VaWqCLtxu6+z+pcXE+6YJCS8MFcQddgkuEH4uW76SpP6iCV6/Meu33
XbJTw/m10zMkCfYcmF+rnVpydhnafPmQr6anN4AKwSFqnaJ6XnBzbpgtrE+dKTAYWLPT3kQHhO9f
li9tJaJYS0qhqNqPOm6Zxwe4CZiXnN0gKW7BdX0ga5qC/2KUKV8eX1xf+aWBklt323EoEg11vbeb
QrntXTIVQWuZgv+e+dkIpLdhlfWosWVweuE6geBHxF1cqwRzB/6fcB0/fLuR62ZQcXUXbR1WINRJ
nqohPJO8jqMISANH+NTa4z/kQhlTWTzYv9Fw25Ju2S7/AW9OhY6ADhUXhZ/NcnlQFq692f42jcke
7ISxb0Ok9dDtYn6vEwIEmox/JKNSsDsiJ009swQG+llexBhCubM4VsEP5sBr+U6giVuBEQMgrvUV
OHSd1Ql6EqchNurpIN2+k9JHRknctH+EfRlcJnfYXKfONPRq487CYgYwZJg8IDJk8HK1y18nfVhZ
JpZ40oRoTz+bdvAyCSvHz/h1jX44pIsBLn5bE0JF7oLmYswhwnpaMFEPc1msHRHT62QGh/A4tzp1
6xxLN0I0fgLFabU1bdtzWVCGfDmLr9lypSdkuy0GmdcY++6kFbA8+He/GhXmUXqgbguk4MqmsVT6
MYtrC+CpWjmadDVY+TUwsSYWzl5m9pVaZ8XYmAbkbhPJNOox1bFr/xHozMXqYIEhqtZq5kCLjbEn
O45a41o4iq3u22fQCsweUa9jWOXGh8EPb9UhPR6jp4AfHWr4A0I3MdhEOlcd4PutGEJxxOOVS1cx
K3S560PqabD9U0p0xkbCxm5Skti0pdsdNnUA3pW6Jrs7JSCHnhGUfRhK9VMDU/019tkY6VT9nqAp
7lzZ+kFSiLuWcrcmQdp8peSoUtNZpYOn2p1OucXg9aQP8zYCZzRgi65zkJEcAN8138/qqG2hPxCM
tQPiNxpxsbc3uZ7/TE8t7yGpR+D2VnwaIi39uo3GRDpD3mS6Vp5M114l3Pg5C6vTR3FGejB9GOtn
Eegy0bQfTGmBp+zMv9gBB81d1ZUC3dGQ8oB2PjslaSa/DmdYl3HVNCM/L4V4+eMVIocO2Mxs94Fz
/BuPj+exA4AqqxwlcieWcNxzTBK1rWbl1MpZoyzzyRDFEYLJ3ry/ArM+olfnmQApz7Dj/CMacxe+
7YUVSXXqb7pU0T6NT9CZdeyrSPdCwlseXH6LfjYEzEJC1DroXqZhrXb/2pQFUssUHA6IKFl6eKtq
NCqLaAMqlBLaWyG4jcz9fG1NzVkAI44zcD8+YyABxfLUO+NxnfA1/j6T9sQs1capPKIXmHe1iPCt
/IPVYbUfEgpQnIvuevP5oU9bBHAr1z+ZZLxlhelW1GS/lT2gBKMvpQlmK+aBhqqGSie9xezLZNrV
HjWjbBoDnUbm2pdMvpQYsqj/9tUgJjsxxKtXlh/+qwJC+uxFNWMXeXA7N7OV+N1RH9c56zR+yW82
Bg45BTKdfrcG3OrRYLektMJ5XINjoAMFr0vk8QfgoeZGK2OPjFpNuNO28SfCVbkSxECR/Nd6ZNwD
Ee+ELP5yZivWTut+kkjZ9MAL3hA6EPbSwknzWxGUyp+hiPPrx56+o8rdpvMpAMeKM1Glzc+Y3TkB
6QvKdc/RKj1jbwVq7DLNDs9DAbUQ7TjD79AQQr8shttSMjyIKYOczPcg1n/2SAu/r1xkkkFliKUt
Mcd6m44ABytIb6wTOyU8k6whG2arqweUacdt2AXotdQ1dkT5OaM8/6Z1MrGFVsOoR4EdqEv0icUb
XQ+5zYh826ZyQOCNXA0R06Hy8biZORvwlypIPCRu+VEzKYujVWeoPa8Kzby7bjr9Y8O6YYmzTfXv
kc7I+SgzaO52AnnIfWgydTHfK5K7ekFamtj4zSiJW/O4qORjntA8RMszGUDXX5Q79FTqt8DUzcas
IT2FfmH2ncMG40l7h+MWdLHgCK30D09yEnaPYmW6qmXAZBwV8DOAPcKERKJKGIBwettG9S35OTjE
uHQQPhBmHre21j9Z510ScsEFPqkTeyRa5n6sgKgRHwBURHDBFCxXj3sx+fSUwX6VDE9Yts5z+rkY
YHBcN2Bgkp1p/G6qNUDP2RVtLA0pwOLDC7NLScsUja9oOe9WZyIjjVHWQ4xUvL1hcGwENSbwNo60
9oJjviw64z3mwdFEaW+7aUroZ68NbcWxUu1TA04ktWQGheqnpQ2boWdaInO0VxWFQAgEANQzmpnc
hsZPTDvgIguMAZGjXDJr9ptHeCmJoR2WUri9FoJnr034NJ8LLOAknJsVYSfZ2I0KfVrr9J15prF8
13QqVneeCjG2c3+PiQU0I0B8ayiHobTh7uMuuqMPyHSXT64Jjv89FbHHItlpCPIfMO6oiTjjde/D
wiWudO5txb6KuOJBl7XzFHuhN7J1G1YumNju8jJ7cC/B1Jx/d4jNWlCDQlA+Gv6wirDKBoFQcW1r
RkCiYmNGxSzI1OTnt1PE51qoWDo/kYgatWQ9vCnEoigpceVAwR2zgRwu6RZUq+lTYSiLSr4XCDr7
3fJIoayLzrXYJyapQ2Zvi20cWD6MYR2xhVpKN+bUIL45au2oO0FCMTginiNZqwrVJ6FSfN5PubyW
ByZLhALqEBu5DSVwwb84362EjRqn12qs/mw0M4wD8KubrMX0qVwA0RGsKuxAVp/DkL3CIS88kAtL
+6584oD1urbbweE6sNU8C6Unr3ZFpULve4q/e9XIzR5Af0xg6JNlB+S3hu+PAQPSPNiumB4sZM7f
mh7ODu7OK8aw95j3ewDv47ksMk1rqjGWGYYPmHLmFpVDU9UzgI+3/DTqMFtYnMltSVZJUHUtq9Nh
vkXY0r2lAnvDpvEBQ1KpP456c58B9CquK3rXI2V5I8E7eBjeZHk7+VQNMn/oVtvhqOitvUTsnj44
pIi37+JGiGgQ1m8sr/2hAfb90DJ6Uj79CmqyaLwccbfUdY6F2t+BMMbAAHU8Fyl/PusBxJ0/YnBf
LuXP6rl3CZPXynYDJG1XZlw/EL9pTewbj4F8Ybk7Yrsval7cayfSgJgBxPZicgeqUBmzCECmAMIJ
mZapI7htrT/z+4/5YcjkqFLNeBkOdWhKz0TiAPeC2J3EZQ82R+usW6qntHYgwqw3/9hLq9qEFoyh
Tx95iQL8ZsugX695EOuwrzzftVgB/I1vNItHHyAy77ZlFciDOeh5kVRf870WGpAKbQXoJYc6NFiG
avW5p8HqBNBiY2VDX5Vl5riyx5HXhsRnbgr73ILw56SdOg1yamP0ra2jDv4uRo4bTZwcpknH+b3U
ddFNDywzzECWYcWrDSCBL3PK8oz7FlmloCR1Yc6T04grRtA15eG4J9ydFFEIoqpcKQt5SxCdAUYP
ro17ZKnCRYPtygY3ZxsIIeelLTeWqYuCZgVaiw7sBVkeFfSMwVZjZNOftC6nzq3xnTGhbF8WGXT8
S7Wkl3yTuRGUiFHTpJJMP7FznhdehFnZm08oQ4dO1S/kFo3ezcL4mF7nhuObMCGAJIia5EeMdzG8
GC1MIhPYVmvZ77UJst+qgHGC1gBhqV/D/CN/V52zyAfhDr+7n+Gdos43SQPJKkoUMTl/xH+aY/br
oL263iq9IUNbDpXpivo/cR1j3y1nttMR6VMUZLewEN/kcpY4ZgAQ751BJ4R2zQGNk17SnOGrL2e+
WhplA47ADLZDD7wEdb7sF/U0AO+UIN5dB41Dnkht1/ludx2NlXuY32j6HnAh9aub/Y8M7pa5wCmf
3uHMr9t9x8qmvA1PuLHIMylEyV5yQp5eiSSd/jllsuaRWxxY/G5JiuWX9+TAzyXQEOvDZze5E2Lt
POV9W4dBvJbiBQNlfGVUnlOU7p5Zs4OrPP/2Pml8fATgDyOpQdDNe/N/qwjVMiQQ0cZZXI+9fcNK
4pRFqsWTcy+wXrFSStTtxc20+VL9kUv7lXhJAqHyHuYkWxOw7xtlINDDbMBujt9RS33RM4zQOHkJ
Ey8Eywqb1WC6A0tumv340YJEEDZOclBGxdnfax3AWV4qPy8EDdzxszSiNxDeThkp5Z7wnd368ybZ
1Vt41d9AwS5X860vy918d1E5arrzuqoSrBwfXWB2eswZy5ZBJvkjgunoc8oJT7g8WkWIo1qcDLbv
VinVtd+uGicykEVoyFGigaM4ovzFsT3biwQQcQj9PbTsr+BU1CznR+LGwv63GdMOLFJq/sHh5tOu
idTXmBOWE6oTTyHl52LVpf8fgTuWMsVReedWn7wPymH1VOaCdRwfG13Ba2y55N/92BfyUwdc1DHu
Q17m2YPHhUSTpG+dAEN/AE7tBezKcj4nB4tIS90nDtTRpGvIF8zfJgTLnFo+U56vcYFKV9qdZEhZ
VCXDJv+IA376uxnyCNFi4d6t8zRTzD0xaeg9WPQOlzv2Judyj7nLmpm5V1923+co+xGI3AKhV4bE
LZW4tO/D9O0q41Nu10kg0T8H4A8atDtMSXTR2aQsJaeT3JCGvB6OswscTlrMqkKt8LQdYORSk/Io
l4xrMUyDJmexrhxIzAk3GWfWpqhxKYUlBIWtDBtRsOHyUj+I4rFAGs9Znv2TPfMifHrQqTl/8aZp
XvHONiP9oHmSBzVlVBOi0OFB+YbdNhvj0OMNurXCYx4nCSsx7bPCcFrIxaRC00TJPqEZESwtuGPE
byoaDzJREG9D9f8n6qgU1a093RyHpN7u3VIKbKrLfeZqkFpLMHmAd9s6LAB1u6SJguToWhEVykEt
paTxv7Wa9hxvdJZY149hX5/bNqaC03SKIaTVXqpCX5vgU9ZQV0ybRGtoxrB6ZpJeOfxwqm2FcIcA
EF9y+8byPsr6Dhz4JPnPP1A6EY/Hlyt4nO2BB+mYAi+6aVsVIfPzodD7aloR8G16N5efHWTj7/Ds
JXPan+cQoNxUK7stBQPjkis/JzK4yrtowXryzlWmFlmnGWFDYxh3RUwlWeSjhiPIzeOB0pzkFeOq
L2wPehe88n0WLkJ6yuz0cTpv73FWm3X0xVowdKNwd411Y01bWCxd0o7MVEiKICVMzZrgC0HSgTSM
hIGnRMPOUK2MYuIpPsBgqtjLNSd/fSWfeydWRQPksJrG7sjun4w21epwEocdYt8bUNiRuVjFtDWE
dDwWuYbFrne4Ohim9/79kIrCzVcU1KN+IzvZGxLtsbP4FTw7GMMpcs8nIoPucSt871SuodZ033Sa
rUg9sjFyi5kmXlFRyCAnznoXbGyCXfBIsSqqnnHwqIX6HwbPUlciER+H3HGSQe1og8wXvP73y3Df
FAitt3CZC9+xrhz46GlrdvVQKskfJ7uk9rO7KugrHKftSvAWxZFDcMHce8hrbnAlr9+jntgWZw1V
HvUliQ7A/BRnfOhhyMyxlgTxeFad4XNsoGOAGz3XqHoAye9DmKwkGMCDhzSMrEdJ/6lwQ3ZgJ7OU
rFQEy/TLIfOn3A3LUi7XWOaWM1dljNs7jjsVTRm7ebEX/c91G0uCnZ1nduRXlFgAYJDROVDqd+C2
YHUR99MpRD2uvaJOicWld8FqLTghhLKFNYFQEcHn0FgJbH1Nanm7sW2FOd5rFkPq8yhe3ZcAWm2f
r3Jf+wESblf94b7AuGGdxLqnxhuvVTOmYKzrLeJUgGoTVI+uHcxEj+7m4RE5g0DG3uASgzH4XdRd
nbB+ZdUt5FhdakQooWi68OPEG8UAm1R4l9gAAE+pm7XG46OlTnkd9u6F9/3SgKQi3N192wm1voa2
E1F/jzsSYe7l/enNYehk7ADiHEXPfRyxKkaKqWr4V0j/AnBodU7pss7Qe9WTG7TZ4nDfUGWR/PDa
/ODXz7HqoqWW/hQRJYGGvX5sVR9FSOZefdWaUybeIqi2E5LHhsXq2mVrmJ9yiQC0r4e8q3jDJBWy
J6xatcGYLE1hNWZX5cquiYgVNI0k0EIFW95PRUTDvm87nTO4tKPm815Z6ztoGlXxKGddScpx/yM8
A9V0x9qfm0HU5QUKsRXfnJJlgG2oHQ62JiiELlAeuGzrzx84kB6D1jrhxqa6QF5X9TthWmuu/Gqe
k+KXdiPnjmeGwAFoHoKm2hlWW2x/zCw+p8hYVXmFPFMyZKSAFC6LNms9yYp3v1JiP4/wB5krV2AN
xXb/OYkFImo0mo4FFZlZDW+Kw7xAJvumpeJif0QGDpn3YCKWRC8JJ75X1r3N+w1igrUlesqCYli4
30rix93Xpmsl9HvIiIDUdFnyrcXZ/K90A2qEKLvb5CswSj0URXhSVhGePLLANjy5XtM4UfTFzuQC
dn9iYjlkqlYR2KCHLL/G7CLeDkYtNnM2RN+TewynMRn5ILCfJgXjLHQVad/cm5v/9erawnlis83h
3UxMVmyfXD78JDux5iEnUCPXzlsI7LYafHvCkpbQuvHKt1eVp2jHEWokyOAOaKKjkik7xfuDyJJS
iBkxQIQk499ZDmAbujJ2JgiNmZ00UDhvm4bOSO+23+bHdcrpCNUZj4f+IK/DGmjxXkGVYVo5R8yb
CwX83Pg4D+g3rSvqtbjk+7mwBACre0Hsb5iH4SzZyKC6zrpg9a+Zq17sKPW8JV471/9q0MuDPGJx
A39dX51RsEHE4zEDQv/y7t6LSJUGs2V2VWo9IK97v85DLpNEsznVMufRwHW2nWYL2wSzdiMVxiwq
1xvZHpEmrX7RhYMH2fFdDmPEBJT+pd+oRx+U40P9c45K6wpg0PkZbl8fEoK/RjvIR7gDyRHDORYj
VLelOhI7j/We1f9XpF+IrsZmauVeZQKGU/We+YAuo6qvrD9kPDjx78c841WfxI9ePnmF3wF9i60J
SmL5JPsJiiZeFJ+z8l/JpeU6kFKU/wxf7j5d6J06QLS4jpCA/YFBb7EMRMg0GETuYlMiWXVNxHSW
zJUwZloR3PNk0lX6S8Bnwk2dqwe68Mg66jnJVOJNJjlXehit9KLBCfu9PfFSoYzMI2D3H5bkTXLT
CuuT3SxL4431Ah+4CTcAgd3oQqp8ufOzGwShsVTy6+Pj0ObteYFY+O+G8DNffGqfcpTYh6pNJspo
S0TspSIwwPKDtMys/TJWaSHkbwvAflm+fU1MPVNlArE/0S7gtHv5wWkFvMIwxmh2vhzTuV/Tp85f
278X82FFHjJ8BmeB+5Ioe7BRu+8T6KpFtkvXbgRy1sqtEZNbZ+lof08bROwrIOs0MskjB3Oi9IR5
Sl+CsqfJJDsV/A2fVHQe4fOpyzSusZrT5UUFhJSv5C/rnUpLab+MVnxHUT6V9+cTOIDMb8OMygU9
Kbvz/HTEaqUxTTcTSUsoAOyWrQvdvm8KdDGHlozn55MBdN5y4lrfTy3FaOIpWe2GgzcfLbR3Xwbk
ylyVO8BhU1pk5MElQzhqXtuVna9rSq6+RbkR0FJR15MAyEdXRl7WmaxORPD4nioxqMTIbJJvEwNq
NrHR6zQ+UcgE6vd4bYd52UrwfM0jsYqeUp2CCYk114xdjvUPc7G+AQnMMDpqSZ8Zx5/Vl2TSsWBQ
DFZIyb1EzKglgxMElrj1vSGLBUMbVrqIoXma1MET73tG8h6SEF8wZzxGdaDpYHO2msl/3pDzNwXO
RC/uEw06Kv0LYzzLuKb1Eh5iZeToygu4w33VSbbiornuDjdXJ2PH60IP0vo3441ojEVdNtDPGmst
30znQZx9h5Cn8piKJMvq0V942b68LPyfRv/T8hCCCJFXHVktx4U6UBzYt7nzps/OHFhcrZVzhZWt
RiC/AvGncBd9EKEk+zERQqPW27E0fq2zJp8nF/YNGmY5XTUqZB47EtJUzgmdKLZsKEF3nlQvsBHR
tvyYLDZ9AVZ/tewZxVutdpXcl89b7NaASZd5VWxDZ8PK+VggZ18OKQ4HuiAyFMJ/rSqvXEYCA2rl
aZdeS858VkJuYBlKiucagQzfKec+ek9WL6aQDEfckFXZq+O3fdVxylHRQ2NrkGdljR+j4T9Hhv0p
xoAg6A/JM33vscTcEmS7EbRGSWN5skOOtAovDb0Ot9xFMDdleD5BxvHvqD2MFyBUGTRsxPu4Oskt
/II+NT2SNIJZ7faD06yxLizIz9nTRkSncbEHrv6U4mGvQkRZbm7AWaigVs+ErHmg0RdR8w8WP6jt
JRYidmytYQU4uaYqRGc9l8z/oTaSW0RwyuRznxWxxnN20COvZpFnju0Sys3Ggvxo1WPiz1ZmxD55
xXFQDSUAXKg4SmoZmNhqdc1k7EM3Gx4/JQKDPS2JN2iEEKdiCYBMXCYNVecgIn5+DN2BbnqHztyu
++7SzUSq6L0J9Jb3CIWJSpUgG5mzy8s0mfJNcbT1HJFEhf7shQtxvmEpRwmt6oPC0KZ6NIWS+Ewn
PCNeBCh3r80zCy/ungpnXrIynM9NiPlodnEU8iB0bkySdSca7sWf0aTUUM3V8MmTk3XUZ85C7StZ
fX1a7WFm1c7EwelhvflrQMt3Thfhvy/OUS7XqOLVWDbgCnUjzCdC+nUD0ncrcfLnLMxrszaBDlR5
W2a/JqJidlngdqJoVnVhS7JDzG0gpJfFTf34M4mmbFTbQw2BCW15QPOsC7XxC3NILl9WJKsJKjEw
+NXlohFv/zXl7RokgzU4AGIH+oZyj/m1+SKdhGgFKw+RzJwC4IeIxSGk2cFrRRiXbr1Unj8uktME
uRedjitHt626EMHypZF0VlAeyunZC77Tj7lmy02sMxwfwW05IDMA4ayBfwlaSa5mEruonwTqbi3S
fS54ruH7oiwWwopYmH2tglbURW7m9Ocs07C8iEdH80lWHJqfZ8ESUC8Z5qFGkLKTDRf168Lac91B
PjpO3mEoH1Ubfhdb6hNDFCG5zcKmjTEHKmEymZgqX+pLOqKWc6Jb1LvsZDV6+0ll5aUZIKXRsMbr
XK8xIvSIHb1djsrcCDdfbpHgcfCG6hgdthsH+gt0HJi/7cvLuB5nnqW78IM6uayvK4dXJ3Vp2xvV
8UozpAnRDYa/4huWd7LEaf858HpGvdP2SKoc646lbSfGa8uJppf4KUfVTPgf3RccGNTIjxDN/QF0
xQFkw3ZlpmltBbN414qEJErX59Ifn0LomTzrP8x3ZZXuohUkG4BiPUt/qgjAewwZcrkO6tJjCPBi
P2b3+PRRK2lg08bVBntJt+ESTn+DUyszXQ/plNOB92SVj+eFzSIPc+bcWL0n/hFyz+PBVArfN+4N
OliIijHu5EJo9QjeNCicECphKcuWuOuxuBLdZFHTEVtgB9xfsOdIMwbC9UX5vBD/qAVcEJY5Nq15
8302mXVTWGKOL5jSf7Z/ws2wYbNSr9wszZHfoVjE3tLU5+f58Yx3rrX6Aoi/yL4tRZ1fj/BNIGyS
CtOV6MFHh8IFt28MVkBrF3c5OVXqla39ogE3NRK8IxNGG5CY6NTmrR15bP7/OTHf6gX0SbJHXHNk
UMRI9NqMCMH5Kpckd8Vc7qMoqLyNiHQf4nagtxoVhxAN0whkxOc9UivdwvqNps4/4b17+XDZbAm3
UygujhKDNkSuFDvTy0tLSJLLb7ofHO1Na2I+b3boJl7+ZAwKsqhkNM8i7EqS7uwElugO0yCDdgLC
RLp8c2BSB5L8SzMU+Xm4WIj+pn81PfzKWt0ZlIoNOgOFHMpZ/jxIMLZogMbLh/aCLYvJXVL//BSh
LOXM2DjDGQV+uFxf4a88B4nC/WM/sFHu6t1fw/5lFQVGi1NR+gcYLFzvhsloSfNHW1i5kP+vhsK8
nu8AJrujVOj8wHQakECha+PHpyI/66PSQW463st1rh6lhScePDQ2DrxB/pvNyAgNQFt4NfvyPVx7
MzL7WpzABiFLzz2Rm8V+imkVZU/hIj0DlH276OtHI6iz3Et2M+sKxxk3ribadi2mikPbvpTgJrt2
+jdsfAJuzrNvgIfLlXiMv/XqpQdvoHlWoynXk/gHd1g6r2GcD6jq6rmIsU6jOrNS8SNGmTJGB54H
COQ8Cmy9h9XcOTohsuLqTm8Mw+YZfnqDcl+VNkb1Ck7rR1Yy2kMTlIUziXhk0iowZiuElIviI6t/
CRnU+Fd6/QVZHZ3SQP6X4R2VOF1lA6aKJd2294xrqwB4p5AvFnihCGXN38GCp05tsfuUhr4UsRiV
UfccJ5FFBy0dlKTtUmekDpfS20UM0gJEek15vC3UYXOQ1MG7p17q84Q5KrA7BjDLgEAFHtJx84jZ
9AWA901g7raD2iJDvlS1Y2R/tW//wHduM7760/OqjfWGoxyAD2R1JWH346o3LGB5IKYI+uJ9xKRD
/zOxzbLmh4AWa9DJqDeAIzHGLzATOMxv167TwukjZC0rglTfZsbGeGoYbMCuBcsDQR2u+je0VpBK
ZUU298731P6zttAZxvamnuAmZLOX/0SN+tSN1QaE7I1xRJsD5ej18tD0oS8/E+fKjkqVBk2ao8Cn
nw+brNlL3vo+CJ+uqx8/8CDobkYEBqJO5NcAc9K20kdjJfIPmxamUCfbS0p1OFaMp3bMArpShWWi
vy7kpWaYvobf9+r98vGyuAVRy7EOhv8HQCmT6sUFxZtB+SsL0Zd5vYJfGMqq2s1QJjcxotX6wPbS
8becOJmtQ4bbWLoIZZ6YxVIjxLZR9JVJvofl/OMj8TcRtwUKBnSQlFXQQniK/P+aGhQ94tSr6CJl
qzrwLh5r6elz/9WGES2VaoiFDs2F0V8/Jn0x7b7daaprQ+iIUO8nAY8r40LspYoTzSkpp9RjYo1Y
c+5zxDyMvpGebWXcsIHErNdSw1aGz7aDHTyBSq96ZSv4KyjBZjF7kBesWaBEIHTmRVIxhcRPFS3q
NFXEsSvAph0ey9VqI+G2Nvvo3e7HR+k9On9gPKP+I3P26EiKvq1P40hsOUwW6D0ucxthJDiROIsV
Rwqn/2dLJfjzCHHyT3NrGYkkq7SfBgpPpiiYJqvcjthnlKnB5eV83n/fIHIUmW6psdjaETeYHzfz
1AJmANwhxkKY3hhVz62GrYMgYvpz6eKgiv2MHnfDh1GRAhJaQ5oXeHLIe5uHxHkkhzh164AZlHUE
9lQ6JW10mLHJmgd6ZCiWTuAPGrz+gETf8vZyWzfxFuqh22D+leqY8Bi3mZDwrkkPZqrq0/m0oYqQ
/ehsZyNvgbIBcLj6aymwn6GHgNkSp4mjqiVuOGtOsBWSBpSA9/J998Xs1pzrJEnkVqLWXVv80Xb2
AUM7h52tmBzQXTT+V/07ede0J+Y7hucmk52/MgPqJkUImfqGQJzHTzQQdmUnv6d7Zc+3f7BnZ0Qs
fbrXyNSDlnFNiOAbC4GvmTglz/6zpfNqU5i7IVXkh9lmYnCfcHrSX8FVX7ky0wF8hMNUIaIFxEbT
6s5mIMn19XeTdVF649MTDbBDrJ/0J3wS4zMOKMayVTdjzT492GGS7BxwkE6zXf5n5erQdnllVfdY
ir7Hj3SC/d6wTHRSJF67Y4m6qxdc1Hyf0bTJTiGXyowutIBW5FYQAWI3zOzm0gowF9eTO6+BiYvn
w/3mnoHeU6wCP4bIC4i3r3QHwS7CKdlpuw8TF8g/V72zPSLmjd88mSbD3kbCqZTQwohHYETVxtP1
5IjeVVltdhvlf4Xt8jhHnyzYR8A7+WO7VoEK8z09DMX7ART0lj1aSd+GEKLaJtY/qdAVPoneKZ/H
NfkmEuZN05HZe9FBaKAYH4lbF0hFoh372EzpYB1NM9XCl+urzc8ieNlivAVuSfDwKMbqavw6ThAa
sxv4gZBI9XxoavbGB9upfOLON6BJWvxGyrdbhz0VXlnZo39tN5mRR4hdFYbqTZSapogGzFAi/bPL
W9ZHBuTcal7J/xyi+ztcKI6hfyXGcLvbhH3ciQ+v5uKtAG/D9Bf7MuO7Eyr/ib9/z9V4dqCj3yBv
lFiMDlbDewTWp0n8hXnkKGGYqdOYnVufDAy4QqLWUZOE0M6Dbp1yFbezP8TNCn6wvb0UXkAqAsyA
5DYizbH2HnB+EViKslVvgNEuqCzIRL1K4sSIGr8TgqmvqUdlSZxKoxY2Kgu83fP+jY5wT99pjJbx
WzQWf9th6RIfMCYxdyVXBLQwlod38qtIaWkZ3w2yIOrrABn43CoSW7OAg+aRec5CxESOIHlwo98r
R2OVTl9qgtakmoc6aEWPhWFX4NvSYUcYixc5D/0HgziMQ/OB8RIXQcs5voHOko1gyVXK2uO26qO0
1ixYozj3U3iv5AN5e6ZqeVLBKfa3uUBv3QWlPVpKJcEVaABDX92CqMbxHxYblqx1wgWIQLtfZI/z
ypAixAYXd1EPpB/WOs9T9ZLM8GCly7wMzn4sUPeZY5G6zGRsXE5aOlV12suAmkbUucnfQZMPwHWO
8PFrzn9MxC8oIh0Y5myppb0eoqdKO0jWCkXPQ9lEMwTWHifiBPwvqOmKCFaaTGyw78Qr+uHT1GQp
uGKLINRdyaCbrWEKpr2yTT4ol4QxqTzpY6f5OHCDlpsacnkBCEJoP3jgc5vVBErLO/u9Qi1L6wmz
+NV99RzXt9yXZ1jZ8Q7U6LuxP6YpV+XMTo7rGis15K4w7k7Mg49EmuntKD4Lx5noVdRLtCwmjRWT
Hp2Pg9/0S0+4+tB0tfB7iTr6O4KVE0mgwCVBKCCW10njPzvwoVLuNB5/EBaXGZ7EqVnsBqYifnAg
sgdsGqU/QtL/Gsiy5q2MyBkhf1Jid8dCr2X1HVT7DDiopWE5yb0ukJ0c3YwqeeKIW8RsKdC+dkU2
+sheAc4RgGBu+SZtXl4pk/XwnWutod95nMqWEj3FOx/nFkT8U77dJZLAByJKFJeUkAFbs7lb+fu5
6TuwBFjG36v3xIe+Du+pfKV+XdUUs83Q7wr9zzAXs2uR5VO+umCeIUV04sO/wLT0BGHhYVQWdimM
X/x4T3dyuS5VLc9h0x09o5/HKjgMKPeF5FR9X0FDwH7OLVUR4Jmq+viNAH/Cyfc4NaBXo3UayPxw
uEGj6oI4waj4puZiVwCywqtQUmFNvp68Pedbicnzoqvbzy5poEPuzYSBZ7Q/BZzFC0+SQ/gzzPMJ
mTFSiI5sfBNAsNN6GfDdM1Qk7oDuspMw2jNpf/xc4tKAT4EaM8xmRyYo3ROJaZR3EYNidLjLXEAm
9HRRG2iBqrFiPZluLmuX6LkNbbnTP4nCHMYqQB8JjIm/EpiBdPK+GI8o+9O6Vv5WLiqNr1CiUqDu
4/PKIEHoa9ldUexrm/hybKpMLrzIH4wE6I9jmRx5ooq2mHqC6oYKAjD9di7U6iVwqf3etjmASEOY
zXzB8HqbZHlEB5XYAUuZnGRPBwXw+eTBqIPKea+DOHvsF+/rxO01IewhYJEnjv7/9Dgc5qGG3Wyw
GYS6JJ7N1jfAIWHV1oxvHA+YqY0tWRSx9GlYZZ72HjQdunYJmB6+cfSHctq09BwbqXzmxdSB0G7S
af5agqodrLr14LvhhHl449951/U07yjP9UKowFQhoPL2vhvKD6XKs/dCHxraazkBXFwCp5CnK+RL
s0W7BTDqwaHxZiczeH46hftpYk+/KzucFsJXauFazjOHIWMRYC6ZcVeZQcVvJp8wHlhDlDvS2VUc
NJ7/cT7wv6dN34ozjBNlBw3ntAeQwoafK5Me8t/yT06AXs9Uu/CbVC9KWnhFy2GKkvCWAM/9XaBr
V3HkOoyRsPSAEzq1yKN3HxCZpI0IMNU/8gFoK8glQd4YXCMrAjA/ey4iGzGhAkbeqO/L3LrZKg86
HRBCV1R9zx/GW+BIIcYByDlXaN0ZI/Mk2fMxql7W8o0agd4gsCVa4ffRcCO4Abrq0VRLdug6x0GU
83MyLnO40hLxJtgB2Yfmd4clL2e3F0tMZ1kSaiSn5+5YS8yuTg18b/cdKF3VKT2we3JbgPmO5x1M
QA7vPXseVjV1SGZjwXIb/NfFgjIN/y3I80mSu6+sna2aCCgNntIhvRpHPZvm/dRj+SXyfVQ63UwB
J/XnQH8BRUqKQRTW0zuz10acVfwfEfMPviuh8Xzd+eE7XNAC1Bf6YA/1C887I0uTREw06GHIKnks
MZhIwzkLewS59SmJNP3PTR5huLv1WiNVd8BeRF2wzUcyGTRDrIlLVmZcOkIRV6KbVtJfB6R3jsbk
PCpKXmRaGOzJoZ4rYx9144ytO1EcMOJ1KGMgbR0APpnY8mGQcDmPQC6LP1Bh8Qy0Eye+AyekO8PF
aumjkTeU+m9wy7d3U2B5dsBPiVgf5CdUaMvpD3SRLMUBh6EAyqqJDWtcSatZJsx+v/NqJqWg7KUU
Z3RsAsvxaOwBW9ck47BAP09EEORo6Oam51H8G5mq76k1gfyfhTNpQ/h+rmvBnbP7n2j9EexGp7u1
LksX8TBxHjTikMKaTXzuOBYE9X012NYQcVKvHrCCPvUJhtuBHKFVq40X0eTndkIB7LF6gXTdqQDH
Tpcjy6j9sxRmjEvxVskwgK4sfD+agWRTN6ty9UqvOP6/RqI6LTekegWBB6prKQUsUU5cYTCNWFfQ
KDlb34vUnKDp7TjTUgOVE6z7jYRTABwwHDKQ9J1UEcTcr75p/DhODPktyCjUuWDmG1gKgjesGvuF
7thqK4nivGAKc82xCD7VjNh5bbWnFnHSERw/3apt2EYya28bFF1/u6gG7nYsDYv2jQLZAihI5hzj
rIwxkHZRJkN7PdKg7WHN5L19IAP/GIK7z6zI4hC2xXDILbdhRxiavMHxxCsTqyMXYBMtNYuD78Dn
jyOwvLrCaeE+bVug1LUi/xwdc+wVhtfAUcEEAxPmEkS/rBAQ8xe+izy5sAruezT6xW5XCDlarGxK
DSCfCdIbJP0pqdygjr2KoH+0P+WUhJEkveE2XoOsfeENSSo+4ktXn2x+dp2LmvV/8bxXBaXrBEBN
W0Ll8n74VDuqT12m0P+o05Qt2BrxsV2KXAKzYhfi6uo5pOYVdpeziz507ii5VFC1n5k6LiZQMiWR
XqcxB8LslmE8o02+JB0y6fL+zVXJATITpV/a1YQjx+/gVddt1t/lvT7usBpvYo8HCKs6ocbOp6uI
TgkXi0O7UK8F7ZCElSkvci8VZXZ+eMhDmc39EFi4XIDrdZ72tzkCFqeLGcAkZ7RthY0Mg134I3PS
wMRGWhEEmZhZNba7deyxT2Xuzu/xqQ0Ca4MMj2GAKTIJnvY9hzeVYFRX2Xxu8f8zucAJMANb//Jn
vYtF3mMx/BNDxUnRNMAb/5fwJjZR4+tn8B/AKFdeDsykMiUw3jqFjAgEbmBhK0+GeUPU6uXfizpK
SQKQP3qdbFXZFmxi6ApLPBw0/c48uSgJnOLM2ybT8lxcGrI8lC1izlKprWEBUNktIYy/yIF/UZ5K
oulrNMGT389cppT6X1YlQTdo/uABtCvoJZ70iBoISwv5fVaucWMAc9/KkqqZhcerG9iCI3O7L7Lz
hfVZkxnTJ5maqCiBaZxf7ndw4Xyl3p/FY6QqrQsPiraP/BZKAufayf6jzwq/1ex4bRUv7cKe5qEX
XLhs9u5BC4XnsP8Ef8Yl+4DDMF04Vx/FpP/Je2ucQh6lWonxnJYYtrbchFMWgoKOj66aknTjetfw
uGuL1ZA0rJ+ABCtMQhMMzWQlnbJ8jQxAaWJK4jfCWyFtiZYmS/C+t8DVRl/My+TKpavosia48XNh
5w/rQBUicENBdeS015RlvbYJw2bsQiGypZaKCkPkQbCs2iXq4gx94h02krCeGN48xCQvccwELR9o
bzCsDHs5ze1JhDF5CiegLYSngbGxM/f8adZLkRzfl4AfujS56izRWH6DpndiVk7VlK/IgIxZwFjb
3aOOW7EDMwtBEgs15fgY8EIoUCs63GpexvpWNl/40q7tLMoPaJNdRGH9X8sEyWZ5tIOcsNiYMgHc
JJfmHzZqgjE0zISYi7yIW1HXuIkMyvaRnGustydpi8UPrWMHCYw9SD8H+sylogX6id0v5H3VEpcs
6P0vUbeibraaJce3WDJY8Mn+j7mOICSBKOXBcBw5NbQyiqB9D9Ap993smVPgTF91TUOwjpPPz2T2
A1vIGBX/+wIb/1IxqNqDdmVLexkzv1yjYT8tK6M8G3E/AiQpyvWDCXuiepb7kAU42/fTk2/SJSMy
8832IVZoKtUADS0CTBPMP5DWTps+CvYfHYozl/VQu/jnzIO9a1Fz0iwpIRMq76xpJ/npseuC5ueU
bZbTSdr6qUTzjTUvIzJo/OxQI8K1ign5Uzvr7KejZe0hCTBWHH4eSt/WypNcBNoMz3ykKEi1EZSR
+zoU1h4vnSZiqXfZDcXCAVh3DB4X+zgdE3O/jIGkcySbZVxdPdEeWrgaD/9L8iACOfgmJWpde7cM
DweH9YHS51ooZUdHBINXEDiuVdsTdGV7I0ELClY6Na2XuQxkEHjGxK22mMFhOirT1fhUVaSua3yK
Ge9va5xjWGeyM917Bh4EzQAlZbQa+vMB4rqtIAAQMiwlZqrPhw7HkNJU1Td/1QbhaVsqk/OSppjv
lCZ+5H7AXfI9Q8sJ+oKzC2Ivm3kfjE6lQnVt6Hq+F/R2OoLkvLUHDVGuI5HMz/7o33P+sg+H1oQ3
eST8wuv5Rm3fX0pm0JwTabGlEbuDmqDliVUdEi1VeRAyU0dohtorH557jGLFfyVjBNzqwIkcTOv4
pbKCHUVBlaw2dIKrR1TNpx2SGnW7ES2WIIuuPCFpB2eae6p7UCgS6zD0IRXUL8Zy87o1eVbWXYby
umoR73+KS2lk0gqzuLHO62YWd7IR1JAsPxKKsAP2pK2W1YGMmqLYdqKNwtNtspapBMkDBkLqjQzN
lZfFZ/s8E+OxRpYoe9hu4zrR0uB7Lq0XC4cVUxOsec3K4mYVPDe1+6asEdAoIQe9bFqvjrHFI3IF
0gHAXw67m0qgG9GO1UMxA09jLDv5gwiUhici4lr2HY68ay+I3/y+400cSVGuZP3HZHUf5/3T2BFO
RJdwDKxLGTzDxzFTWjBnB1QypZvUV3vKubKzKDmuw4HxedT+yizg6yKme+5C2yw6OmIJRxBbkwc5
n5f527rXZayk5Dq8G4qYnKr6qmhLaS25n4mcLipFGxHu3qr8QShNeP2COyXhdjAKhThfZ9jTD218
yXUD3+8C2sa3AhQmuegR50h9IqYLPvnOWyHt4nQLbRDrY0skwwmvKaM84VJ+eQnpalQqqUMGCyb3
w9hAbcUFI9rNw0zWHg5Sh69EITTetvFV+BOeOjTE//iCw9qrpHcpD9mHN3eVJ+j2Rj1Rr1FVPHLB
MzHr+LGDX0rM5Kj2tDqDDUNfU1uOP8bafWu8HPcLNsn9FL9mbPFAp2T1Sc8wedFTaFZ3h1006n9H
sBXHzUeSa8anMzSv3NlESdr3t+9Of4p35fTrOfTyxRxrV/M6Bg7nwB/bnHyjqdNhz4J1plcYmhns
COArlqz/4lUlT93wtY7Mmwvy5aDSFYDEuHso4lTK6f9KHXxmYCOIB4jJ0+HvCtxcsCRDJBDx4KeW
PkRgMkx49hPD+6y/0GDG9OpQo4nhpxVxLIK8Gut3qcDymiLj628vM5xNbNTYh/lLIHq7dJqwNOcT
RQuN7ogZQ96kOKlHX+S9/oB4dCi7oYlMhDpA+POTSsovLUF/gxF21NGnyhT/zdXPDAEEQbFq0bw5
zDMP1KjrajGPQC5RXLQhlEozwwD5vYEYahIozabyqMdS5ywIsALsgqkiSKTkPP0xtLt8PVLcxb4H
ImCbNEhBYquWQzzJPx3BK22CKad28//1n7Q80iSrzMRpuY+tJd1i9NcPwLLJXX4wWDCEIrn7ENIA
GxbZyIx4plbjUHXQWbTUPQVxAClfnt4/RPTBBL8pF58lmr/1wIYA/16718kms4LW17lvfeCbx/XS
WhNlisBGUWERotWESruWRcx4ml+b8FTIfjijgnoGj4Dwesjc+Tfqah5eoJe+sQyzJ9ux/d8hJ0eb
2fkf+Mw9tFUR10lhVqzhyU6eDNpj/Cg2wDz5OOTlN+89rDb67su+yQ/KkfWRoYcHRWooXMZa23B3
eLzLq2xJCsXkd2gqS12UmYm1aByYbkNiXyP4hXpuhtQrsEiIvu4V9bFeHNshPjJXyxCe/XxfzkuN
MEgWzopXDwfdtl+JshXVddOVzCBv3u79hO6NYlhpCeQALna4pV0wJFpGIs8XL359JN/a9bpeE3Lc
XcD6zg6v0hk+kTGt4p8nE6+G61ZaqSPYUi4bhOY4ObIzBjtFA2jVU1bLTr0P1i94TFtNFzYxvPtl
efp1ZDmMMgECogc1RO0MrY4VXHxqc7hU0CxceOzOg686wnmM98QEEmieIiDGBlT08L1Kim+ubQnR
6c0nI4wP6aAjE3PewqJLHG46w/VifuFmgk1muP6egXMpP6nxFdepYaFF8HXkFrAMWmgX/3f7l68Y
TJ2ZLOH9x2ABDhAwfEvj159WQlpWrL+Q8iUnHjEQZU6FfP3A/JoIikXx26IqOJpeaGlezqvtWofa
mBXZHFUbm7ygKLrlddHOjnpTv/bV8FSOgT264mgmkNWzFM4J6AuoHIUY5MdOd4Dj4JIez16gAjX+
IhYAebvKQJhX/Ns5IqCiqPV3orG+kVqI+ZUrZ5orqx+icDIY5Q6k2HA9jdoeF5Qc7ngRM5SEsuMb
o11F/SXyELfH4fv3GEpYaJJl5OHoGjBgxTTkogZMy2JvLeJ1JgKVlYkl9hpKnqND/LzcN1HMlPQK
u+WnRcW4Nj9HIT+2d+H1v2M4MYsVsLYNi6rE+/Tq8XjXmZKjXOB3wbsD66GcKdHZJ8MRDGlleEg0
PAG8d5pWKGE/Ga2UTmFiqRsjFKdMbVHufVJ2QNvBl/SZkXs0GwORvMnB4Rj/MgGEu5U0fRaWtMeq
AdTS8s6AH+prXgkcgYinCXDYyho5cZqmsBfT+++U8nHtr7NLFMpmiEdamxOiIo/FSggJTPHbGZ8V
D6Abs6ac+u0OYn4Md/GHeJXScJy07QPCOlcW0qJoLJyLAuNw8sgcf2MFREM4nVaZoIJab8DzSUEL
1nOQUnB63WcdtlFRfXIvpXPe8WT0mCRIx6q7W9qKHjGElTr0YPjYjk89x1W5Bss8rk4xI2Ftj1u9
ONPOdlpSLpHcUW8AkUJKen2ypZubRk5u5hStKTM3RAOMpc6gMXBDz+7SWmHBqlPl4kGjsq+cPDDQ
Ci9HAil8HmjWk7AFpqAwiZhGfLEWEFM1oLQj18AeAlX46yj9lBPlefFCSFBuDtzUhqQrHvzPF5Up
1flsivayereNXOn6jeMpfJIZUsEkWGAXB1r2pF1Y7R5nBXRVb4MwF0m1ow956PXMfIm0u/F5sKwP
NjhPz+LCf6OgN0HfYWK7gZbhf8gctz4g9mVlhMiskCkpdl7G3XI9umivGPrM6F0x4gcvUVfPuH9m
qwkfiAdqEG2MuqDMgo3qdgdGXrDaynZgXJYNRUFVHh9TTvM/U5Q/kg1zPnnqInr8x64I8CfRHwew
rG32DOrXFiMBXmgqGaHNGphSlXqgP3jeDWMpGSGC6FzpS5H0qKBKkqUrFodQ9DVEM7g3fF6oSEfM
kP9bNmvRMrt3sKuAQTxYx3mFMiaOQcEz/cX0r7GWoDKDM6H39OQavj9x8hIUK6wY5FaPFWcyZ379
IFBj/JHe6osWWms4blm05Na5CSDwEn4xREjC7zFI9HT2Ih7xbYA9yF4ZwSbF4cREjEXtZNhapTbp
/htBbBthB/Djf5OleZ/ErvHaY5LYEsfRjAYoXAMo+qZv5ri/9shSA1XyCOoYMNG8JMVtXWYse/VD
qD2NNYxfg816vADI5P+cGYIQ2U5gUX5+jZgHVdb+OrTt9NQVgx9K+ofW4JH5TMGfejXSAoBr3Qvv
l7oBZ7ji7BkCbTyAqVJXYujhr3XIx2A5SRrEpFGAinSfImjTZYlLO6PlNPsTJ/fFHVWoJkeIjbqp
EJrG4VfejEorY80V0N0pZEdx6x7maA5G0utyk9nFjR9LKiRgT/67LgNCyKO5FiC1+idGLUFA2Wpr
LyiKLlnpOtXXyxtT6FcGoEbpup5Azv7vUQinV8hEkeFbqe8fY+yGahR/xSCGpdBuiTo1RqRu2O6k
opqW9t+XoyZnAxsQbfSqffCtRclP/zl0KMtwWnz1XHvpYkqiStLAsaqo0XggrRumtthIuqET/ZA7
9m0SSIxYybTPmyLcbsY0Y+TXUUr3JIW/YwzHBBmE2G908gU2EsqcOJ3wMOl3q0L83m0omdrBKmTN
ln2Wjs8KT3FZZbA9fneK76dS4qxkmJwm+emMktiJQN4E197ioRtC4TRMf3W8CzWGBXcoRZpsT7mD
l/r2dlOTRDwiCVkzS5JJB4RQ40jOsisY7sHNDOfKOSiqAsb+0wYfj9niVRd9uU5X0EV40K4vP19S
fFr+eYHj7wATjS4qhJS98HclfOtyTX0x1JTQlBsnMCySWm29w5bcitnNT2P8jLDVzfgo3BS39O8p
5v0m+SMPyryIqbUrFdpWdoSrKbafByfgYFIL0wR/7qMv8t621hhb9WBqaAeyiC/2qsHpwrMwx9fH
B9tuRWbmEKwzbdjwqPgPkRCrxhZaf89Qw+Zlmti7kPmRCDZ05r4n5SRoGYxiJ8uygyLf2ERkIVLZ
Wd0EUVtk3AMxyJv+DxiKAOPeG63w1BZZecfkr/0PS2r6EHVLq7ISaxu2HTZ8g4+jveGlns4Beu3+
rhRpd629LVCRfSBatqheYYlBOwvcDK10fdrYpnF8SgID7pHW4Q+UgHPN/69WNC7sRAWLmAZkIDXJ
/I22RrgdQ6u4T6gpMUf3JAxYRPS3JbgR62mSTDdxzfM9NBRl8OO+kKKV0n2JeDgfgaa8ABMj+XBy
8LwyYsUByJ6T5Ce5kpBDbUJ7lGQGJMoIdTlpFTf2ZdxrKqx+IBDPWX7Az2AeCryAyRo97/uO7hw2
LISUfjw9Up6PsMdZqJbNb0sTpEQIb2NvwnADhDsxBNwpu09iovQqA/v3Tf6+aaBScmpvXrlKxpfG
0h55+LGjQ+8b5OwVHanXDU0b/vx/EyhWCVe2ch2P62/fkESnPw1SRup76MmRQxWaHTW+h89WnZne
70mb2PNzLrBbSZdFwwW3O77Py+3C7f2zwCGk9vMgT8HRoPCCPhZdzvofqmYyqpjm9sZBox+8KMnY
MIC1lix8AS+WnsuTz8wOuNCwoeXJ2skE3bZ7hDlSicwt5M30Y8ZpTAJV9bavO0S+MCgjqAKKCQB7
obBRWBztNYwYDWCq4HNLKR38mLrE3TvmQo/3ORgg//7kEVwk1Ezbo80Z3eqeM0TaaBC+vt5IVJdq
XI1YsjFxEVNey9igqheF7b04y/xqL1HF9ucRWM7C6jyMMlP10Lca4ODak244KhaTEuuRggmo3D8K
X4qqFOPvTL8Z7Jf+EcSy+wfWIZOxj/ZLBHnfUDRUmnSfIhw+JDHGPE1WMIz6bAyEKa2Wm5a5ll9w
tZKVJs14To/yvGSQS5vWLwpi7hq7+brR6eJb9ObSHVqduG8WzeWgYpkQFbVl3ZdKC/vMyXtHpeZe
YoBGIlUboyZQ7YTjBdZsuF3PiX1ApOZArONkUl+PXIQYGy9u80oY9VguV+6tLYIMhpZWAb591X+r
eR5+bl25xzFFUylar8dFVTvun7BkJNFqiil/cWbu6V+PCz20Yr9hnHhzeKc7PlLofTsaS21LAhYc
1zUdGx3oLdxlgAO/cuuPYaURytNkHSh16szRHs7GNkWVvjI6D1SiEk+i5vHvPVx3sAmAuYlJ9Qmr
iHHMqWXunN7BGHkbnRfu0t7nixwdvrpLFKb3cC9awri/xkGt7lLaau7x8YVszV8MNkfCq2RSxzA2
Yi7zHjGWHiSNfy5kmebRy6sSb8QuEhlkzucfMpOROHItd1+DLz9q8WuCvJiMJFtMhkLMuGVgCQom
6KqySadH7twqi+UXIh260s7/ncRlok0A3m2ACT2Ie1lnSdq1lUv5uki/hELeJ+/1XaOUsVpuhFU1
ULghXhzNPJfBXHaSfi0Pn8HNm1m8xpF949NWOcTawKpkbYZvjXRkZxG7+zlYHnNVADEjhtapO1Z0
s/f6fB1z9XuWV0mni5ZheF71GDR3Q9yZ1yGoYCA2fBbFsmZWi6XL9rqWWiB6dV9Y9WQRqqy0jNIq
bnW+i4JBFauNOh3T8qC3iIi3SDpB0QhMWt2RRy3liqszqjBNw6+JIs0pPzBT8+R9rgpYQb5iPab/
Nh1rWlRNY92Gj55WrKkFDtl7ANTZGxAwg8VnVrmfe97Iw/ScATHUdEikbfiMHpfgeH67RAFR8OI2
vqu9jJVC9fw+z+pcfDdoYAIhViz8PnA9phbK1gL4a9cs3UifQ6CDFCXHu4t/zuog+m4hGFa3XXIg
7DEktdZtdjQDT2Z0ljAWROfB8ZJDdo0V44trx/pjCa/n65ApntwUqfOpxgpULAELQ1FiOgMDqBYn
h5AreTNOGU/WeDi8kKQJ5TbA97Vw8zrlTzEbHo+ISpyrxVCILNEop4SxcD/uVyXWPo7tYZAKD/Yt
VbW3mqRWFCXXRoy810oi+LA+NvzSF0LPPa7aj1vIWG36pm+fhR793aSI0rrgma8pc/mv1YKIFqVx
suoHHIAk8fTMHsxW8gzWGJs9KPRLazjwfIS/cKGCSb6SRcszTKbZemUX5nqa2QOXpFBpoXQMKvIz
we4btcrWfFJtzsfw9LjpsUYL7z1dssMSwj5GKVBcRzULMipcydoNjhysZ7xWymSelEwsXd7iaeFh
q4rfPHFDHPEYeqmwTf11N1s/jfqcDErJ7zdHRw74yryrMCE5VpMivTMI8WHcQif7K36xHbSB6ULW
9RADm4nudEohQw7RXqSr+DDSiloo/Q4httqdOiVvWwkHY73vCV1v5dHGmB3xqdpBMIfTg0BXoC5t
A1k8f77KWAFA0IX2cl+qody5kJjsM66zPg6CKNNYIHDQN2z5wUnwaDEDt+pA01a2aMtqcYDe39jP
vA5p7Kx2XhK+GaVTvf/9YbOgeoXA3bkomRxxYobVKmqBojQOhQr+XMqQVYYwAKHw+LkjaCf84Yqz
Ghqx7paoJzy+Tt1DzsGFPscgyLtm3XRd1j8MvokqTi5ctPkT9KKutJERhC9Hsquq1Az4akZPYGWy
4yDX8jkWDpgnxypBfF7uY79is+b1oagN+L5KnldE2yEchZ0GFr+T9ZcoRrQeEjEs0iKmdiiaTMPP
QgBQhV2qQ7Cp449mO/PBbvWUElZxkAaToBIbZSh7aD+dehL+x36IFOg5NWp4JqdD/r7VjEOHgYow
AVJ19/mOTgxbbgRrQmQ1SCDP2dceZJOiWItELu1ju89HDyZEgWOSLk7oRw0G7sNMhDJPe9D2CjCz
wwtXsfF2JnAiJaYGy6WXCW19c3+0Mf32lO5mNjb06woWyevz87/EviMbWd10sPAyibfEYzCxOy+W
TODngtJtStk++lfuShmccnBJsTeVPV6XC85NLmYIi5XBRGqLqKHMEUCUsMYxf849IaZ5d1B/yVFT
tV8I3SfjvfTWyGXirZi7aDkMmOQiT8JU8/UiY1xAsuf4+RCl3LDkccFfJpeGLvpuM0E2ETcWdBQn
I5P7GXTKEUt0y76iWSFRdiUUofd27bxP1PTPUo24Fkp4an/S7lOZNe/FrvF+9Scc1BRe2loPuIKh
DqiwU08bKhmo7x/rSdSNFJgdCFMQvTQ6d83z4rjxAx8cY8EQ1wycBD7tmK1EAmk6GSDOSOd8tDlr
R2ICgmhLkOsmBBOrxB6FuMDUdCzV61gq2433luViQq/QEytIlDk57YqU/xzOKUxccEc3pIMM5EKr
Ldky4ZLRPdIUhPSX+5DOGL3lMsGWCm43MVUGZCmyFCRIH1pnI0MKbTIk9OjjYNkbnZZh/PNW10KK
h8JqVkaAjJZTClGvo78FDmketbyKN21UqacRQCBRBr9QxEEYUUDUeGgmqltIYcwWTc7jJzewXhPC
J7SXlLumMjwrNTPlvgh43GRXJjk8Im5/x4lqCXnk0Ce/DJieo5MhcEM4MmCEwotztN/chFX8aNV5
itZNK1I+/gzc/JBb/UXjnTk3h2vYrg9OHWq408LGU3FfR8mRM4COi9glOp6W1z5AmZ8J5qZ1Yzru
TlauHc2sZBDaSX/RA1X3w6OVnXDNP48ydgLZ68bEeYhOKKzr+YQjaGkfFIil6omOY64R89kNFqfL
+Q6wqPF+QYZFXERiK561O6jK5KBVNqJH5i2gr3NIUx8kbH02/7tsJpH1HHtuDsujv/fnpO3s+FnX
GgUkz6baiXehiqmnupLIwJ7+bK1AXSuqq/1k/jZySqKZ3soWUIoZVvDru3is0xs1OR3PMuHtH24z
HGD0hYSHK+L0z/Y0ylcOpWv5uyB/wq3SAs2b/9KlxV6uwYs5s1sjyzVi22YdTJ+xWm72NPf7zFBZ
7TE61aXc6HtDHn8G6od8/mLJWUUJz/ZE97bv/Xx2U7UVIc9upgJCSmqNZ2OsYiQb2rkcUNHVDo5v
6DAie2JebFL8rDu4W70tfbA//EEk4zVIqNFdvRaQ7tVD178c/8Bu/dCc8dU8zaYD++Ka32d7rgau
U1tqSP4ILAAxTJ0JhQ58lOcPegYYrynZ+5JQeIRIL/PCF0QkwUby8DwUWJ1cIaEShj+46JkyOA0O
HjRG10Q1eQbL7ggfchP59wnTSYtPEnZPXPhA+UvchNINnEjmIsQjPBWzaJuuJJx1s5FBQSDJYknV
3AhqbNG+1fFPsvZuF7OW0hHnP0MG0wzXot38gp0+AtCk1kRtiuguxHwHETiB47AzwyMTsSXMLXlq
P3xEA+dUWNEiCnJOuZTYKkCYxJk3X7mP6ltw72KgWnx+JfGskahQ07OvESLwTkI1OjBQ8r142gza
HPM5XPeqbldTwPukJL9KbupQSxs/NYLKA7mvkPRHAEqRUA4cCPxXsjNxDtefWT4eYjWribmCi4IE
+WccknqpQjX1s9zpnrjSN/BNZSgfuppl+WcLfc6ziWyqERHora2mI0FMTcDyYesAc1fjD8aq/gB3
9KLVQA1ScknjvJPFMTkQTwnhItaj2zlmWsAPLQsGBx80sTbLF9/WAoNKNgQ1qKiCvtk6UcPdcp2M
Wki7dJEWPOl6KPaMPgNW0shkNkYKc+swrV74gDaIcJGIr7aGro/HNNzNaV6I2DIGSFzF9hxIym25
xiblnKSfOGzJRxORcpcSpiojT/hHmwkHvm676jW2JVWA6wE0507Cf/hqr57ptoLsUye0ypxKNdBV
MUinzrjYIEGbZJmxjJmYEyeZcXck5E3VgoEx9p2QGQa5KUuFNNfDnuhfmfHHkA85WvcxiFWARIc1
XrbgzAoqvVwEUf4q1qNWYGC/qUmkg6V2lToN/sDTqzl8NB+4HOq3irUhE1V4K9DIDSDg7J7nPp7U
ilui4t6v5JwqqWdjgAe7WthWFHSs8UFWOVIMCPfwKOglpfPRLcI5VL8cIv2CoKI3dkofL0b37epJ
Wb1N0cDb2DRbk8Wv6NwfktWLz/5VSjg/VkcBBSBrg5fzuoCjiQSZhIUy15zBXiNYnVKNTIZC6AFy
cXafL38lxn+ydFusol/Y2BUZjqvbDVF14pBljKdVboBqgOSuumcy5ikuWXtySGqz9zbUPJB/nNOT
5iMvJ4cp+Z4d4iw/g2lIR8/ZTnwNjsLQ0MfMmLEEFy/cjj389wX4677pSJ4jg29fUDYtALO5crdR
w8jTADFD23NBTQh/iZ+z7xmoRsk/V2SyfeZtKzWLa7l0j4ae+XEo+aH4eqE6JAxMosKgNSchGhqi
p58OQF6O2G3+XnM7NPY0AmfkxyxXH62DNCvSQUU75LH7iIMsli0nkjZh2CpTBDshFKFwTFfj3m0T
zHnXD8tyV5+zKD8oYiNOwLAz4sjvskeXi9tDg315o5+rPrMHCgpA/9q3gEgzjjJjTKlFp7kkJ3yF
gb9t1Ny7QSal9w1w1v0E7nk41wG0onQ8uYASo/clYfRk1mTkobXEHZVHKaaRsLtoCjZ3NpkhL70/
Z1ZaIjVqWnAqrEG2aeEpYttu+bmh3OaOicJT/wZIUN2TYrhJhECc/PVOMQXP2NpjK4RX9IBMZhpk
8J2rndKUW3XSeMNtkJT1WQr8N571TjLEcmN0xM0LBUvThTxkgi+sJm15gcg+csZtp1BB/PvBFbnb
rd/HzKjhu5T4rA+iF0RI1IIc4I45QGPKuKxptc2mSXTlalEZdvTL6chQOF1UPGhKiAP4BINd21aU
iS/nGbdhXl3AYpfrZ0GbE4u/zELq/Igssy7Kss4OaG2loECZ9wcTAfXlFWqf0GxZNrLCmBvX8dBS
ZsM8CaR63Gw4GciT9j2IsNzXrW98NfzCfTKDOh1EUFtu38kfsFJFrbniStOoA9E6xp6+kOnGgNJT
l+21mh8aCxE/q3abdJ1cgR3+0wqLQud+HA1maZygH/OQHe87wAZLgDe2eyXF+frW5l7FbgnZNWUU
yNRVCoZb+pEbWG6rimEEwzo/rHfuLQSLQN9nMdLD7wUfVmM/dFSeOviCL4Qa7Jd2Gt271GDG/pJD
pRUxRXMHR9AvS94BN0MHZ9l+w2OIzqbUuq70Y6VrnkI5hhAj+9L1TQ0MXizo0jnq0e1qSSX4RTfM
0+IoKTT+9Bt0NPA4UDc73JRz/+p09hOILMjKpL1HfO/FTpdWIb2/sp6lObPQjDarpUuUAqamUBpv
DtOKsmjUDaqWALdUHLXiD2i4o9iisaN5PaGWuK3+fMWlI6C3KjtE2j/zmfRh84NAhzl4bt+6iKYh
4DmOHiP2ZGqNuDfYtNiGUKJUjgz/JPnsE9mJb1eNf1zQi3DJE7e2CQPh35Q4WWGIm9XQ2YfsoM5V
wnZ00IFAImPxv0bsbG7Ofc9jz7QeVv7kgo+1cDtq/bK40vceIDOeUiHkB+3cXmBsbiivTh3XDeAL
j77kR0Hrh2LqFrzxxTBY7w3+GOApzrMKYXGxOCJ50zXWgFfvEVgkQE5gRv6LurwFb/7b2m50E8Ir
S0aIV6gOVIwEVtp+GnO7ZpgO7nhsXEuRqPNiLDpEE0cuDc19ZjpqbpZDL+mi2SYL11rChVAerT6K
tc3bBAba75Ye93JAHCUMcG7UEwwhVvKDW9UXV+0PmBLxnkQXeJH1NDtynkgflVVhMPzduIPmaCrX
bsERmspj0e3Uevcwg24/SiN82eYLZAWOibaaEj5kpWv0mFsi/NAZ7Z2gY2Ijs3DFi6I1XUQapu9J
ttTAdgzs8D/8kelq/6SxkOmZ/pvlF/srX3dsNvBRjIo7tT7mQFvqovCNIkysSxbsxoNG3wXW3inf
vPixiPv7XbG13ofEcXegoPRsiCkmue9ELQ2OkJVYUsh2iKs8v0l0z4l8l+ImrRYy7jDQ3K87A+Rq
Rypw08o2TvsHCR7Zsm3QMRGxWii566/tOYjhcMBn0MrEhqCDCIFcwabRgai0ATojLv5E0VKT0jny
nL7YvmMuDLIt8ijLylG0x7DQGzc9xqlveT+YA7jPMUHm3u50SOBAhHnXzhgTg+B49otmPsy78r87
lgnEtY9fgwdgjg+bejkqqyOjR2kCcSmYXLR0rXg/aIXPST5B0CsR9kqA/1X17qQ9CKHFHOHpNJRa
ZUjUPGdeBG8OuUuJm615+VXgz79UrINBmYBaQORRiyFOuSTjM9XH4e8/PdOqCxr/mjSfquPizEk/
UktoncglqrSwdlcigsSj73g52rVY7V379Fg7KA2klN+CJwK9fOugKCSmnzvnS3MTSEfNdJw851NS
oGABZmdF6MUBHyIp5SsMpw+8tgTP1IjCgweMMsSsX7gF3cwl27Ku5Fs5mHVQqglHmdcZjsD3rLqM
7Hs7yyZy1oE5NFLmAAlvC248DUMSYNvdim63rZIjeEiTNV8pdbJKiOYIayTiMCW+Blla6+BNLjbo
eoc8Q5POcm3LPV7vLbK5vFiAY598a2JcNa4cAQVRufQyI1H7B3+VGD8Xwm8swf2P7oXfBcdh/V+7
2P5SdxtjLefZi+4EOuHui15XgW4CyD9KH+5XaJSpAmjdeF5oDDmgVHXk9rGAxhYfREKIRc92FRoy
SAq5Bn/Z/PiVWi6hKL0zEhWVwOheM/d6pkX4/6eAsvqMviB5vqkMvGWgPTEnHyGciaWuZPXNEVht
DHnsnNIdQ8UrO6N0d4nQgSBaZU9ogl9YPTj/smjHYfQNc4+ZFVo2e6tNt7UKpqEoy9WPXVj3+yvE
UL4BkQOBndlpjCJoYVs8KxqKRlJuwsO6Q6vZ9gOBeup8qqxgy4L+nyDv57uMVayhOEx131FdHgag
6iJrLkSuIBppc3VQ9jXcczBUSEu/hc/5UHSDNmiViWo6lXTCNDzoHaEcvhFxo2NebgNPNf2YGmDb
iMCgK21+aVPd0NdmXmNCVTUlGSY1h7kd+UoHf8ys1JD082RrIFO00OJ2K+1pdofYys/YDG9gVDyc
FTxnl11HsWDD6M6/FTYbOHFgXGrfg5yyEc/LPs4MB7TBDL9AmzeknEEPW3VMGpUu9lm3ywgDJTU8
igXO+oIgpOffsFn32Hsea71/Pnkm6EaAYFyaAgPT9kR+RJRd3w3rcwLEkZffxWF5HGmi0PLLpIjJ
3PugvM+F9p4mzltEtJHQZEwzPMJLZh2v6PjwpkmxtjdzdiOPwZ16iwQF6kQFK7fMq3wLqkpD4pX9
BqRbqC9MEKdvJsADwa3z3cUYZnDQkB9URclvdblxS/tP5wZlDF4n5wkkrdM7XWYhtZFhE11Gjg4G
a/VREGLL+ITFWQhZm0oBZOFfTEM6b3aMACg/J4CKAxW1FipG28wkjB8kUFmuRR18899CxorPru3S
JQK5PYDrotZpauxZhBRacGwNwqulGLYGE3Qow3KlUZOrYCVZyeUwD02rMzkW0RWUTwgOmpgHb89N
V2xsxlLoBL/QwrPdTf89nmS78aHWFGUlpkr++SzNrPPuYWMn1I0WdYwv0sKrZVn6QNhvLcQCFX7U
BGEi4jvpCtpdUdVjyTsPl0Evq2nLZfts4IpKL1wIlqcbSLMDoBMpV513kt+WkYPFV9vVx/cDuXM6
d3B+4qcI/UdSqKEh2wEFIFDd3MPRVBY6zS1S3sIb2Xp5cdFoLCNVnnn6qWsyewQV/lnjtRgEmZaX
wpdJS17VVm4IlXxFfl4UWZ3HpU2/lQCCEakZWqwaMLL08/ODebnKQqqV9gouQ77EmVmUCikiUaYd
LLClovw0DRwRCFoiyYIxYewB8ix01Kd47NvhYKIFSP44ZUpYtPTA6lOwj4w53mGKZFvzLR1+TIw/
k2Q3ptLdN0sd0v21uT0yehKmFtROjraudOD4HDCQFIGzJgk9h5piEFGwcJIXnHYOD1uFyvSR3jX0
Nrtsxl4BqBalpmyn/DhKaI1QyReGlrPpHl8tM6IYqhIavzCLFr0B1vLWFpGhKI/egr+sdLoxCUHv
LolYoBfYVbDBbLjlYM4a7FqHRAg7sz7P8DhXmo0nstCRnOyUEkkXMVuOT5A7JDBLOdG4dRolAvy5
9/g47Xp6Kmd6jYANJojxP+bBKobZg+kTveAwLuPHlFoKW+jQA8k5+/LghR3CvqRXHyuOG9QfaX84
nGxc57xGyQyXgvdUoAetfH6Or0uhGHB2VnnoSLPXBSl6DnxzjEAHoPJi+FTnt3CzYZl0kZk0WqgZ
u+zD1ASa0rMxu56uSWuZrvgT5SF2hMTgeA8nCWrkm1RVq+PLcXrJPxDBplOLW+O721HLlH6T12gk
XjTELCybLZ85qCCoD0WMVxzRYZU5LNQatnSJja6S6Ud/f24Wh6m4r+a02Jmo8a+rZuMQ2t6nom0n
ei9fq/onT2PIeYg2bi6gHNmMwRONSpcLoehUSMW2ysCgwiQwgVHs6/G1vwwCBjIKtVidoT6rS7Y5
h/q74nSTECdv+2MOqChgKVIw3dl86UMfkl2CwmIN98UJNx7/xPY1kRTFE9FP4iLytQfYmIP0eYhn
ku+aicRHdh27l7SyF8ezpw/+xl9wZRjsso8xiDQwFeveUhXv/Ij8mSXbmd07N05Mbhu95K2f8Qpv
SEmwS8tYKD9x1YgZX3l1BnJIoisZHI4PV7iMahLVhQj42RNHOBoU9dkMoa4wQuo/q+Xoco4dg3vz
sY78bdYPyRbAQ4wD3DfPf3fgzFxKbodprzWW4NyHWV3JzGVI4QoB+0csxOiOhZRTD1/rlPetJqkM
x35lwl6V19FXPSnTmOqsL1le7ss+cmS1lkT4Spduw2sI4pXC094kZ3ORiR0A01GAp/4Uo5DlDgVI
HqvjOGpKRCTfCKWRQjkiJyFHYnLdtUkGsXZsJds8+HCg6dNJrh7Xg4P7WwrnDE3/dXTmeEqz9nYa
rgv7AYlm9tjYvTrLQvWzBUQ8JDUVS0hRxkKo2A/ZYRjDUp8wpjcchUl/9tNQ/lLgLykPBmoM77cu
QDFGOtEdrQwWWhpWD4HED00ktdofP0V7hC18W1XpiIc+TBUucaRd0ciOUD71nSHsrBsBbrL97ISI
agCEM0WLI+DD8+YR69ZY5pRWski205udVrWjKIR6B0SYJZBHlkuVfjH7Iy/LaZrn7Y8nAF6JMf7X
HlZWSO5iq9sm/BW9egoiuIk+5LeLDEIoq8lIRIPDxYt5UDUma1ifyWtOhonmt9r2z7oVV0xkdYZ3
xyJYL/SZsNMmnljuM/L7+QkTcsgvnoVdut0wS/dgw3lkESh2WCgTAvHy0Lhn03v8D14P4Tt+3Jax
zAB76bVtImKm3S0/14bxD6vIPUXR0XpxjY2U9DzWno3Cw87MduX4Zi+9JwzCkzUThQ111+uGnHVO
4Noj8sU0zkIUz3IsF56TqYLqt3tqr0j4ddk3AVR3mIr07XEl2z82GctwIK1P6Lkw3qSrMNKhmpsE
0h02JkoTQhFi8P9OBhZ13xTokVbcYT7vx2pUFVRrgkg+P2002PsHIUD+YYkUuUMhXIk+Y5MSGplM
Y+uXviWh7uUa4niLD6/YgeFFLA0SdQcujL9OFxCl6b9Fc1cCliiQ8BKru907J6HWpQNbIv8OIb6r
OVsqXMVHDKCcbst+6ZK/act5hU8c8FvTAWVsvnVD1yFHVAHGESLfU80jhpEPWWMPkTPMsAaCSE4V
asWY0+CbetnRI+Zn+JIjRJ8Jl/Z99Ul94cpkPK9CmxyEFeZKf1AfARBaEUkliVI5h+JTVHsMh+Yr
SfkuB96kiEc6NvkJNFInU5wP5ALbMYLKDv2otWOaNU4EONxlBWR6nTxUlLPrtb0EDZ2yiXOlvHoR
VZb2s74Q+fNdRvL+RIimo2jcbrwhmDovPjFPmZtIBhoTr5n2ZTdOqr9GDrDZL0I7H4zEjyyJ/7MR
FwXDf9wIyzQA8TigoLbT6dkr5sUE9czAJp8ce+YPdhUW+h/MUpc7bkTGyvQ6DLGxbqUi26TvX1wM
ta5UTWikmhTpvYLET0csYKPwcM4VBZsQ3DcVs3YWXv991YZc9hqenpuw1eP7nJ89hA9j6/b9Q+tY
4M5hAQ2i5xPXP+i4iUekk+GdFigrclRRJTAdR7QdzXetwqRfAr8yYJSTmiCENJFPZyYCAbX5547L
50Ag/Vp1RLXe6MXX0QIWU3TkUGg38N4VcmkJa1cIT6/eoyIZ3npSzxWw6RVzzrHEkccH5bWjj5mw
I2emMvd9fHqaD0ULEQyOTJHtr1kAM1eyo3RSlHkCH3bN5qx9XrDd3Gd3NRcyRvu+iYkSNYBiHG6W
9YC1HIiSs9eTE4IuoDgN+PncJ2YoHHFtNT/O78QxGW5OYNWbZV9jmTXAsAUlghFeonziexFqDfEJ
4f0cOmIcps5LCRW3jUnnsN+e6HANKFp3+rgQX0rXMwiXLVBVwQSK7Tb6Jnp2rX+AaLmR+9ydKzzl
8KkgdQ82PBbkVgadF8Mpo2fBEXi9/pCmgk/MgLxnawbRtRLJOV97lJZc5NJ3EkfQ2eRXy1iyfLE5
lgqduw+BYUUT+yGT0S3RUUdpo2sXBNihuaDa67r41EIldljJfGCc/NHvFmhuh4XMZbVLm4ThZ0Fc
0te5YTrLQB1/20wifUGid546k68tPWn0GVjn9DgL61Ku6JtFdk71IEFGe3jSL9vHAUWBOjGuk5Eh
Q5J0JseNWsdsw04YRBK8hOPP57HAJpQOqv0A4qo1Enb7WnPHl6aPPoJLhqHhkaPC0r6mQwIuDjY+
zNakRrT9H6rWVmbS5KOc8HdhJtNwp1Yz+lywMuhcS1K15Vk5otfvaamYuqw8ULWFS93fZNlEhfA7
qsDo1f/ihxvbjO1ZNYLJWqkQcwDXLrjun/WpGUDMKVRFAS6rkuHKc783NAA238W6TrqyTxPv0xZI
ymzpuZ41QuSDD8tf4WIoWqU9uPpHoYXi/W9WxNv7FW2v0XXlSX/Ov7A464nONMN0TA/IGPKuNkq0
3V/M46e9v4V41sdB3rsn5x5Alp7BrjoBEbGMYf9ZQzWoGZ/His+kOjBbXCxWuqa3p/fZTkQVPkfj
5rxMEqtAkkB0RFMcutLkXzk/CFdZ3Acyb8LDfBhAX2vDa49Riid6eBapXRNGEzZEdmZp7W08IxJN
hZRwSljhT1wYCkF8aYtG3TA0WXf8pxmGyZUbX6fcJ0ipS+JCJpp2EqBd+xXNzIsc1+HypOtCIz3z
D+L4Q08uRnv06Aely61q/LdlLjVAy3si6fEpApd60nfVFp7Oc8VjIZRmca25nNb6sIyP06YFo3Rq
ihz8TsFvtv/bEjZxZ4FRAZMPnAEp/5dBR5/PDyK246t1LoONN5t4F7APTy+dHq7UVUMgtRwQFFez
Bi05YrXok+bFpehRR5fzGjrRQUBGl9tHoZjBl80XwhWxWcLCPRVuJm2xRsGtC1dpJKXigVrravOj
ykpH8kcfmOvxSnOO29XH8K0ay/pMxk9XrBXjYru6oyX14c0YDYY1nUPZWMUKITMQPETQO/TTK2xr
8SLuP11lmafysj/VeJ394ZsQWd9Jx4qSBDJkBNzegweQmtYKQd/h/xjEBWv2BdcmCKbTTmy5EcU2
ZBsNuyL/cragGIPzZZLLipdY/YL2bGy377bodK8LWp7Y2e1uh9mwSy/dQOXJ52TLUUyeJ/U0pb0c
4LnPXPLNtblh3WV4EoGxFaHE78sMJgkoH2dlCR0Xvu3Gb5lEySoCmATlkJKqcmIqcS4NEuz+nSDE
BX00OpUfc7/xSlPEtO8YBWzd7wVoTKNq5ZmtMTspjHh5HaU2R522zhEpnbxJ6aYz9MOPCzx4y2Tr
bG3ckBjfmCEUq/284KElXVtkF+xthovBBkrjPEa2QI4xRPAFD3bCN9N9fPgksn29qA1qJRJPKPCN
Ew/tABKjBWMiBMF5qFhoYDpxpfyeR+2aDsGoCOXjWsgrEIiRjHbr+mLwVLt4PEdElMR7UsTwjNYm
9Rs0DY+jiIXxqwvucdoJTwIsUb+aEkjc5RfgX01wRdHx2uWJQfwm/09JznTd5rC7+H7uZNo6vxW1
cykpDlVp5nC+VwFZ08+s3k/RZDMwQDG0cgrhunk4fWMi15+TDHtcCN2F8gZHjEBJxkPzuD+UudU4
4AsTS3nkytcGOUHz8xGjhnagUPfg15KSCLEheoyoUQKjj/x8QCgsYCPIou1Zq0gMq2v9DbKZQYQF
gO1ABx2qmJSxneWPsAoueZnQHmAUEpuDr8QeVyVgGpo0bqJEVCzKeYW9F5UVZyePU6H5BooC3BXf
hE3eW6laV41v+H56hZXXGhSYpNmxD1zAbt8XfHZ0Bjy7ZjH3XB07eWA63BcuNtqvAORozkVUwzb/
hupG2ag8Vgo+gVsov/3fqc3VzbOwgXY7w5TIeGxznvkXrDTNMeBSCLsYhtDkMRCeGujWIX8hczEZ
CMXFCSoPQEqRFd4Ldq3e+fWb/A4BMrPMpBsMKWsh7Ot2bx8wfsrgniue+jQAqovI9weR/Ynehsao
fgf3lOtw8R+Q9nrY3a7lM8GsyMny4rDqBODaRdbc+yJvVYf2DzxtzjlStD4uoCRhCsQA5MZKxOQo
bvnPpwtiyLpQfI6kgAQP/O48WhMue/ThSr2Bj46GkSfe/tpY90iWlKwt8Jie71tddnroDfrEZisv
FukiwAmyrnR4JrK9HrZjfj7iHZxoEPPS6v+lwwD6YdAv/cjYWzutsFev3RBzN4lRJZSK2GDJvEjS
KVpZWHNXp5h6fXk7HVDA9OTYiSMSCqWWA7AYWEM6AIDpekciYgo3HQJbL9iAwwJjPY0zgIUXSgW4
618AZyGbVeXMvwjZ/ohTEjnRz0e8rvXYRs23q6G5X1Px+RPDvxQqv7u6dqFyfhUb6l5MKTCO6Jlu
oYURNB7otLnO8mAeyptVRUamoV6sQaTxVNCshHCipNbwBf+s/btZw4E84aMHGmPMzxHCmpat6bfP
gGwI7gwOd/6OlhGfwYzAKN0I21o35FXTjFBZGE2hppFguH9sEuqRXdg+Y5E7jHUoabUvhRV/PUrj
6K1WUt6FID9JVy5sDyEiZ+ksaGOjYO1/25lz3ZEky4OjChJNRWB4wyJLEj+9NQtkZePEheVCIaAa
6Jgb6w3qgwap4MJVP+55t+ei9pnjefsY61bppBsY7Han/f/KQ1J83244EdCgQJSDvSsWLeaC6sCb
76piPiANnGk1+UOjjPFk/yxICdT6EgapXunjg4v/hlra7Ws1N4Z+Vu+eQ+B5onY4YZ0P1pA+aitm
TEv+7ojxIpPuohC2SxS2IlhCiZpjucIz/oMQuyC6mv6DHTZAgDlY3cQMH3p6Y544mvTPMphQNzBG
VnG/6qjEk4C6eSWtn9b5tDbMpJztuyeOZblwDS/oYWg51IVsYsJ0U78iVQyoM62lVo2szaayL6vr
J5cL1zz4VJxWfI6CIQhHRDkadEtr6XFK6sj3AdYxvnC5MLus92efhFsKIYd9JA0vP8Ca7T/lq7FK
knffIJv5uDgTxaIvGJt6zWLLiW8aPP/wtUirnyiM4LQ2In0nP6ix/aZeB8NMb6QG4Avj+jlupdB5
cK/j/MVIEp4IgwUEROtO+yBUkdew+XDBYsepWRMKCUUq5ahXNiegGD3I0zwE4K4O6vvmp+2e/daU
4E8YM+8+a9Y7Jt9HE9EETah/9/ws/+WyPqREYsr4rE8A3zSeeUdq+iffvIXDdTmCsSYLpmW6NLur
YxORqJL5TKIC+aS0+DVe+oroLnj3BGhTj243a8gepqwRZeCEJomgtk0U7dUjxjyucdgcesCb8FFv
m9rf9GBT2om2gnUu4iZlz3gTbYv12dhvP0RZIkxsfUtuaLbYPcSIxs7hQfsY9CykF9ECIePMVV27
Fslq+OacQalu3xaSf/lbTRw8Kas99lWoeiv3vZM3QvTLOy6i6JDw36tiJ0JBighJB7Y1Fc70qd8V
T22GJNfd6jDfvUwheVT4lM74D6sMADh9jpl8gLgQ5DaYlyC8Jka/SduyLJ/HLsDE6OmQ7uAOC9DW
hhf5d73+6Wxgole0+O34DgMK3aN8MzWt9XTA7fodtAkNRkFtGJsqFQGXWw4GAtNR+6qqsVEBkB5W
TFdds4ra0/hzHybXDohi0Qo2u0iqOdPIKfMZ363W6kcSTcuCEYeh7sv/fxXrRaNrbZ5lji1gU5JT
ohY0UzZu+6zhDtA23Ot1g7/3u9VRAAwu5RkHiXD6PSgEXeP92SjnysVmUTsW0U0iwCdgi8+etRMb
W5twcswd6F/kfLawX+E8QTn0xSjh5xXLEq3qVZgiWE2/CrHkZNCCt4/Yfv8igP6B2XEDBnqpP5tJ
Iv3VEVqsrftMUZY5CZmpo7nz7FF8VwAOpEWUt4UWupCpu9POeKHs6EapmIS+NpDciJ5OsaZT7c6Y
TY8tDEmUxGIxD5Q0pgPkiHMjXBVU01PvIuQubt3qm3xnhUG7+Pp3he+OmsVnWDeofZCLRkGy5mTm
XxLWskS4TvSB6e7I7Bp+TnzJw2br3iDKPGZLp53lrTK0O0DNl03qpKrylWlsCYC7Ah4TQxsullwf
E2C3fJ8Pd6Z0+ut7M7ZyAzW//3R43KFlgJtdXED/eBnlFkGCVduqGaFi4rgdhz8K1+r0VapNBK1v
TlDMGJg8swz8H+xeAyNqHTpchj9p9H9F+GME65f1kzitSiqloPLuyW5c2L5f66vSaRpeTnweLWF2
M6wWQ795NP9QqSdOomGy2O7mKR16ZvMta71iHqRcnhbGHIVSBvRRDI1JglXyXrpnSGyC6VYY4gqn
RBdU2JmHUNX4qwunO6NX3OZObylA6S3HQ4WgNmFZtEHhyVxgSnU5TFH6BnOrUsUk9zv9O7zOPV0d
ZB4p6svbvezOQo4L032bwwO5gyNpmRPyAYaACczdO3MCcImww7kB+TcvJXYOY3L18BMs0vUAcrti
5bjuppFiGGgQvBkqjn/ahiPJ9q9t7lEhfX7Kmv2G3KxY7q7dJdXil66Ha+VCam+vEarKxvv8Jw5E
J88OYo6yeqWDr/SRomMPGKICCK9OnctttHcmyXEEKBhaLxSw7UIBMc+xAB/e8DE/cCS+nZT4ZfLb
fSVvXtu8w4pngnl1z3pKk6/FK38Vj5qtXe45IG1MdP+H6WVbsfn786Fqqk/a5V49P2P1enXE0Pwi
BA0DuTjdNHoVlobZ/7N1FvPhQx0XqtX9UJbUQEhG0BjXIGtCtXHX4O6lPJX8llqGbvK8QjlpNJeB
P4SZex0Nq4dcRTRkMOGzOwGxKy2HY4kFMf0GVg6Ktft3l0UeAJGFYfsltMS1//fxKj9A/B8pHn3r
C0wPAwJnpKyaO9RgkQ4xV8PdNdD5uuBzhsCB9Nn3HidAvok1zN+CNi/aQtZndgpifmFfz6wK4CmZ
UrJVkw0kfXlalrnL39MGFQUwzp69MYVcBVEBEhn2/K9Hz0IgPi8aiCfVPYhdWD0lEHc5namp1Sv8
SnJ8uDsw2oKH3v0MFMYTvcE6zy/JXsaR8MBRwbLgTvG4AglwesAmjv7plVlJLY0oyHld+MvPcCaI
LjXFVW8AAqAh0Pg6NXjHdtEzcrfxthgzu36wNSviZ+iRaz4FinI5jVo3yGE3RF6l5RhYjb2dHkXy
tOQCOvhJo1oZ8591ZrMEzjvUdEyx/jRjjwJJF44dCV1w7ejvzqVfHkpm1gNHAQaZl3CrHp4DBXwS
f0CVjteIFKcSVamnuxyLhP0w/NcF1GYRF01+LzUH6hySAc+aHtGfKNhC0kwqR8LOFERgtWEeV00l
6Cj02tKhTf/mcjDVovKCDUvNqqOyslV++X0RIzk/XaoffCEh77unGebnZmC8cz/QqNGRhFVjNWR1
QABK8IALOk9YBnuVWMOw11V6UeXLL8VEYBI5xQr7nFTLhZl93VHqCO76AbkBxmLWYXs1d098W5Xy
Oe2W+X1gLlMI2ZMEsAr9eq7UhhLNmH8Yxox+Cv+F0Y03CbKfApv+dbjvbWPOV+XPBcqhtAv+iLoe
PZS8BwPs1Jd4YWOL31cGsy7uteiM6udhxv1phwq+cfdqumeBZPwHmWdKSV3QnaawsVy8BePQNeVf
Ny/kFZ0yZb0jMoGqv3a7vQFPiC2+1+MNxO5Xm29cJxZoP8b0JjUo2evmlfA3P2d9zch9wk0h7lDv
yPFNvopjPDml2KJFrhC+TOjG4yI/AINMpnLpXOEwvci3K+6/tKeaQXLFfxFxjQBoqf5yZYhswu1o
GLwYdNe+z25m5sqxO22NUTHGK538l96XpnKXY11iW29OxIF0KbQ38ViIr4Ol3Et/eyw9c/XTzvCa
D40olROGhZFnPLNrvLa2XRo7w90kf777Au6gq9xSlVguPwzL54OQlbALCc7a1RmlJyyRAZlMSrbC
L8HyTeZ7hrtziTCWuuOyV4IOA45yB8IzWSyzbaGwDhdo9bwtuB22E1J2fUs8DiriqzOIN9PIMlM3
Xn0GCKw1Lg6KQ+iXBAICCQHBIQgrzOSXiFd3jlIFmUhxIdsn6eLkAJdzt+8XQNKV+MrHK01hz+Tb
cvX4PWZZIAVB5LhiqM12vX85FixcbWCY4xN2XKzhy5E42ij/Ge7k2wxE8SL5ga+njt5mavoKUxwu
hgPhO33HjDvwuICPP7fTYIwM9tqPVFgjfMzm+CNMFkJK89jZpzqftdmlA9Y7Oxdee6T8DmAO7zdk
Lcd3619x9EmR1PUbXndDWxuGceVAvVaWzzFo+kqk3QeXqal+WQvoh3tHmIZKLQuQ9u3QtsurJkJV
XWRwP7WzPpuD3x+TRijy8u6rYT9+lzrmXpxI5RT+Zkk0tODOXv26qUGkrsj0p1XShkh3+sofqi20
mZPvyGk1EvqyBIym4TvViPJGjVaHMenDTeDT/MKvbn4kj70Ia27C9TzVEeFbr3B54ANJdgPyFFlq
ksZ89fsxHxuufMVQqeHIwqK88lZ4T5Unjesi7HT1rKjoNI/j5thhh9GMgypemPjvoMNKw1U5hfTd
1Oxm46Hxg6VlmvY3VLQmRlTARb5RTgTOWrKtsP3zF36O2Uf9ZRx/ZogNISpbGr+gRZGQc0to1y3u
ufWwjECyfM14IOokVR6heUpaVYBsaMTZF8tX40xY5niYyjF3V/n2E61H7azk7YA52ShwZfcZ5Jph
yrul844TgbxaS0kjLUF87RHyHybEvVxgZyBOYbFuF05M0Xb2RqQmc+KnyejylzNZnUoMi/6gNX8C
2zBF+ab+9NtfsTjx2dvMAcenGgIDKyc4CsjYt/iIWDXbj2dYiEJj/V05BmZFbz+WI+5uWskUz/ZB
HYgX6Wr7aK35pWG5Wnvy8vsXZm4gidukh6bY7ye/T6ZOxumRKAczPu9j/VO+qb9RCKiPsnFZ2Ld8
tG+xviofR/cGse3u46i56DlxzLSEbEbFXOhzZWZbc5rqBjZ7nuPaHnJT2xs5bU5G/X6mWhSTUPWw
fti+LzMYhgO+k7EUfEOj4J8QLUBBsxvwxCycUd9vcIkaAN3eH8HRtOw0L31PMHQoTEg10EZbDJ4X
Agr8l57WoVJmA+gaCdtDgBS8GX55NLJpjojWcmxq25vAd/SpgXmiEyGp6mQUJ1Wzx5ndP0m0Z3O6
tUw27ltColRMV3Vmn+6rRBi9iZb18tS9ZbF/3O2MwAWNIZagRuq7quEwcJy5mICSp2Szg3iL9nQm
/yub9orGKxpuTZM/ewhY7e5wIGcdxh6SN1y8FfbSB2jpGq28Gi7PWQRVeH2S8ZBi9xn18Zs5Q37O
AjKK/9+toq1cAlsnWn74zqhLr42To0gFciYVwmVjjBcLHwsUR7yLjV9WhZKJvQemm8f22Ex4cw23
rmrEY/CSV+VR58zKYgqJnYQH/rWwTq9mTdyw1d3/YmJaep/OGJdGOGxw07LN7a+UIDCvrHDMmwKK
h07Qg88uAPiP4c5je+XUfOJQm1kC67OFtGuT4HT3Ftqa9RjodC2Py8HKDIM6ZWqh20Om1QaNX1E+
fGmC6syksin2XWJOA+3eH3+aYf5+irI9SToVuWx2rMn4nf8lcX3L+5r1CJXE8QET0G2lBZw/kmKE
zXTSe1Cwym2XUMlHr64r8ZXsrMB+rWEKHIyzuKT9VQM+omGk+xcdmahnrX1fHNgg+aSARrF0lJFQ
0kPASTX94PJBTQwQiB5e9yvpVGhpkg4XR/hx42834yr4aRiRi9MIUePey93Gs+w4riJMVK5ZlPBZ
0d/AjI642LU6SMNWH42zroDgENPM5N7TaLhC+zbkl1pOJvAUyCmq1Bp2WvgYtuSWecGX1ltfU2jm
fS7EPaFGNritDVS1P/KVruyOpzzlIiSGqyT1zJUUh51dXVjI3wAVvMyKZ+YsubPwEmWCWtwgcgKP
s1gb0PhSVqdHbzKqnXmws8EUN/MQxBroYP8+a8tWvDF5TqRL+sEcjii/l7rcRO7v7g9YinACwTf0
XKv4Az2+Iq4eAG6/Kyi1G4aMvEO9gKGsXyOZKZIGNOYVT3NJB1jrhtNVHml3OMDN6Ne50Esz3Sxk
CkDd5DTx0TfZ03x2y4wtuG7Qg/a6lgrCN2Ce/TrhVMQvEfByLGcGAZOl/H8f8JnB0MaP90jsyzOQ
gxZ7CvRjQf1/7gLxxI7nuVF7+YBLbDhIXDcPc4zlY9UTA3oCzP5uQ98JIUd1J5T9qpL0bLo47WN5
KdD308V1VoQd7AjAF36c0FD6trWQt5StWtqkiD1wnwU38yvvV8hNaxYWqLo+RDdbv4JP2NMXiXZu
CFBoA0NJ9bmtBcWLUL5iHwdW5srJ3enIDOMUz7wDrg7+o1FBjJlzUTX+CG+gOBOImRf9AZzXRzyP
xpOfSfV/GnegHr216EeG3TJKkeaK7vpfIz64uSAbZ0ueNUqNuUKGlEWbNND0vyi/RpvL+LN0hA60
ghhtVZPkHtDWzJ2lhjOnv0ZID5n5OshZ/7lLrz7wpzjmK2TRnbTePYEhboO5QgRP2nccTJpYIwfF
sO8UB7zavT9G/YidtbUCFMjHv+k4RVoJur+bAUpq1BxFTMZ5rIv3G82o6GWfQfJvhQzyM2CsmOZE
PMGi0i8bJiO/Fa6t7xP4iMimWSj0gfld8xMgkemHejaXMjSfWEWGIwpCySMtU458WtsbaA3H7XTu
Aq6uDXHp+vh7rzjv61E7gDn5Fh1Qr342F+PYFkKK3UEBrUquiAv3nsscXAj2YdvF9XEtuJZ5u6m9
vQNtfYmNHfNLNrWlH7//NwwJrsRkvcoWtQW/+oKsIxYYNqcIIciBnmrVhSjfQe3j+SbOD3+EsPvQ
OkoXes71wGC8V6uachBnmvKXKU3U0nPteYHsM6oW+7dQmyp2BHIqQRGZx3CZRdz2p+hXee3XJ6np
XZ29VefFFNMhjUS29vMNaNFG4XA2aKR9iUIOu/UW6ViHC8a1Wy8SfetTsuYd1xhf3zi+d/AOQnDf
2f8Z667GLFRztkQaOoP+bv+Pzew7BfNQk7Ai5MWl4RUHlj5Oo3jUIKB5EX2sOgnx/abjgIyMMSlt
PlYljmnDMYnid5588UXxUYDBBzusfQ3NtcQUrv2juIa+Cz1YusQFXgEdTXoT/HOaqIsc69G4uIIC
1a9qhUo8FWzbU8Zrx2FhIIL51LNhWLrBotOld96o864/F41h/glOH94pus/3VTJIsPL/XPh/J/4b
ulSlAzm/Ie3YzRI9AETgJKVPCKDER1ZH75+aL9CdIVYu0RCefk6iqwo3Cs08hUjnaXfdh61guhD0
uEvNQxZ3uJie/JNXD2tRHgq1XiDwATr+gR3zam3lBmve+5zQ87Y0OJkKpSH/Q6Hb6ww6BtA67oTY
pKh7XX+zOw8u6l2r5uJjw7dtYI2cLGjFa3MxjPegNqIA64Atc3wUfPlGo0p6bNoD0fTINtNcnGB+
TNOO2WGua7WhrDIVpoJS9QFjnW6ae9WMQy20ZRA9nJDTRIEl44QqWvXnWRvveZAJ2B2i2nGwnQNc
bg3iOJestQ0FJLU5IrOvFJJM13BB/w2F4yWHLWWgg7Tz2ARsReJeBDPXRmsfkGSCxgaCV/Fixxdy
cgAblbO6zUNRt6wEwJT6V39ihupXG9pbUliGuHMgS5wlXs3zlGa2aaYRXLrmzps313Da2ncOommJ
oBF+tHq/jqjych37eyzBcGDUvjSKSYO1dH+wLQMTlx5akYoJvRZboQR8bycs3CCfqO0pEuexqRQS
mBpUAzEfU7hrMDzww4lSdMeBXfGEhgZVm5Vi4BX9/+gMQhbNRNJ3jsggwPoAQ2uLmgOoyYLeAakg
33tXYdcLvypmznJAev3l4H4gpn+rjfcHgTwHJCTfFavv25Doiia9DlMljUiAodL6INBpVDNkmOnN
faGGL7vgMImqVbayfagFXTW7rxP2MyyhR6mCsORdJIU0Uhm15272uW4IDoWQR+aGO3bh+QJJI5xw
YOMT3r+8v3y0NHheipEWH2nyDIa9hykr8nq6Ue71IQJJQCZb/UTcrvye3LkUPGc5cGhAFpIkfDHv
1/Sc4nSbXVrgcsSlhnXhAnSZBb4v5CafTxU5R9KLKqCfmuT03Re54+YOcbnL7z2svx92c1eoH5Ga
yn08eIDaC+Ib/FXEx0NyOjGQHe5l3aEhCWq2lLf94de9IDqduBkbLvz0vFVTjgnYK8rvA957NCMf
6ARB3vD9GguxH2pN8Rwun2uqkR5sp5bH3Qh7xBuIHC5K1JuSzQegy+ezvJqVNiStHo8QMaeirlHY
SVbfPjbFzWyw+13hubdmdeJwXNoAvs4lEAx3IRnWQ/UbYklBgpnQ68HPIH29jCAdu2+i0vAwiUr2
c5jc1gsLMGC17SguFWJRwgm8EvLmkw5/pksvXrFUqyhI1xsnDIiEYwhPuTfroV62GYobsFaauu8G
JqVYZgfPh8vu5FevVSafwdX5/0MfnP7SOpD8jrOBgUaZHI60hyG3/T9N22X4/XyaD0KAowk/HN1u
FBl8/NUWguwf23wyEjGPQ1RXFMzd8d9GQTwxJ+KbthcSpbzdJWrWFj4W1RT4HHTkSYHuenKT6hAs
98375/7JTAo0Ew/VGS8YwIemSxyKF9koeTcv4v7j6VSbGm6F//AqYyFyfChD/QJC/ShwpZ5HJTFK
D2J263Im4HHegZzhMhs6xqNJ9pTrb/i5bBlUdEq1yK/AgNM8p2PJmOphRDgrudrnmXN7i0vsqHid
LQITRTUJNoZMO7t5TP9DqZ8T0FGZSMLsLtwO7uP9b4uf+OMubHoBu2UKHuJh/h9XSwPTMjAvjooo
6frtjKC8Nku8zkxSMbF2xp7NOcxReb6UiJi0r8PqVtjQO4WNfDlnfxFpnqjzQNO9JXw/6cnh+BkN
VhSS1ypjg75sbW9+17HFQA8kcbgxCrdhn37B0Y4LbX5hHwWw3b4NyK2n1DpF/O4KeA6UFNuGQ4wF
xCJPZarq2hAMYSCxb4JgFZdtcKwQbxKaSa8cpIhHTgB0jF8psoPPvsuiHxt0trXCGM/tjp58s+w2
bsTlUn5CSgYzQpbbUSFS2ujSO2w16ToWIG7+6lrvXgxQ/G2m1GDoN0eUdJkwG7c57DJognjl7TQG
iSteOtTL5IQ8M1Vo5YfSVaSb6F6sgXSjA1EgyoNQb+F+Q7vlP4j38aWxQd0uoMSA0rTjYG167lOV
CYT+pVMcTQo8vlxulwk6ae0mXreigMbh8MEYUbKgaHA68mSQoG1oOdtFMMR6gLZYhe1kVIoRtZeS
xVMSrk6gB5U597+7zSqrIzgi76hy+MuHsSttrjhdiIc2z93FErMhK9nLaOGXFTCXFSTjgbbfFiMg
RfPO4rRQqHDbHT5CU/jO0/Zo8kAxAjVZQomi1rQ2odDJXwgwDBeD6NR7rGHwrln7uNMiQm5fM35B
DLJ+9crXewluOzdDUOxvR6nWLf0qWVTZCNIIKq13XITLFsWWe2awU+xt/pKDunG5wTbkNCC7xb6d
mMUzw1uQV+t63ORTfRjVqQ07870vJnbSuv37VNMoBeeXXPneDXGiDiLonTMhtywDuLGRoc1CN/jT
nvBfxqmXRMeZpZpXbH9S983LFAjGvV/jZo9phbpFcAdTpaIBZBABs+WnECHsRcfwlGtXtkRqAM/Z
a3qCuSUViYafb0eZzODc1bEreauZtQM8Q32/mIp2h36S0hyFpW+Hu6mSgMWwr5CJOU85H6SXtxcO
0AeRNeza1m163HAj/joPIMCG7qpjwbdjOp+BMu8ez8WOgoSilyvm7cq0odwhZILTqR50EsRqMCf+
EoyuklVlgKNS3LoV95tSKHHLjyQqihgZlz7rnvKYzitr5SWZom652UDtibqPs/ZfoHU5Wa/Rwf1p
li4dhznBgP9sVLEqWtnXkgoXAwavda9AqI44WO7/T2Lj/CY4a+dUwBqCLDOrz9QsqLsnhjyz1psv
G0GJnExnP7+Ua1CvNerklv1GR6ElFe3aKA3eXTs3anQ5iJHuPnZ0G7Nwp6YuIVhus/jXvExqNzED
xekNnNRDeJUXTivBVS9z8I//0TBOIU1Z9j157CDKcDaf77m3eB5sN7h31XpZoRTXfqtmAHEfvv7j
pmtzEUO35IA3nhxDkRxo25hh2gCFEuK4rKlaccsmIgsfI4+J/o47GkEEZtl9IuDtikN1G3GVS1K2
kpJuB0xFvsZNAYZwSH/IhKZruaGqTDVOURxlniR/lMXoCdhYqNBD5UmGmWFalRcgKxNl4dnrcUNk
X8/k5rHPZ02ziiGeAO633jqFimQdctyNysAAotyJ/3RoFd1jiYmHxO1rQqaXv/dT+ZKvQKrRWPcr
A1atrIpIMgvygkYq2jNs+/wlh8FP08oENv5IxS4jCqwLO85mSbY0UGU713xuvzFUdNhsdMdkv2R8
8/wciPHOtfRHLhdxT5kLa2KqSjQ9cPkIU+LsRybLe+KeuWqof/9MCqGk5n9Yq7b6SaE56dQQr2zU
jq1hkHTsNNmeN/GPxHnEXqbh5QpNqVXbVT7r2ZnUltGljl/2gbNp+zHWg81JK9Fhb2LEZ2j6P3nm
xZ9GFoBDAW+03NkRe3Z6VnQ7JmLmtODqhcrQC7o+SxzlJGWdVOakChJ02Unrwd4xjTRzdX4Or58Z
Z3a8Jgxs8hxRkmN8m1dEKzhFTIs712EpD5zJfsgGHykIsFu0HHadTtXo1S+iqZveQ2q/dI3LoFEK
RXo5uFXFFhuwVVprCUdQ43xKFYZHThoBemTBeJsia+giHkyTCs8Nb4NBaFEgg9EdRl0XQIPGZNwX
vtY7WwEOr+IBkmRYW4M1T053dalhmUDa8W21CmzuD7HT4jjggmKUoBawQsEjL8pLwOlk+eLUl6o3
45lzwcGgIk4cioqOL3f+6V5aW1d1FiixpqcDFABNEubn7iKhA6awYies3MFAjOMYU70wU0kBwEWZ
v2Xnp+GlvpeVtf1gedOlxyQIa37RDmEFdBjKtDdgHzhbDXfbHFSPlsOUgdKdfVO/+b3CfMY6Vn1s
nJcy0EE3m34HQnC6O1/9lq4zLe2F+Uvqo5WWbE15cbY6mDEhjIisTKWvF/hPPlf2ynH861Tva8ee
4xlVimAmTtivu2GxZwzSRBRvoDZs+4WEKAa8wmFHUGNEW4tLp2yiVCgK6jO9lW7ASaoAhkNMITFG
zncdGamaGGLoFJZef/FHTzxHwsDc4/+QBJ0hl3OPg6RFe/lsR0FZpqK0CV9GyINvhRMMPc4fjWb1
nFgvNuJIeQo47+aMKz7w7H+4dY8YWqqMmWxs5JwwmlQ7Mtl8Gzp3iBRKYVkFeqIjb0iCiP0rajS9
EShuWuqK05HKhyRnZIZCq9+HzbIzX32YAx8liVQOBHXG03qdkjZmzwALQ4B2fLojXUaFnOABRDaB
PvkqHdaHHyAATVxAApNeOZ7CtF7IMgIST3FGODB3AnnWTra4I3Pj/CbNPE7BYwIDPt+kZvwG5NDw
o+9vncu97s6JZWBQ40Ozvi9K01ba7nPLaLTGZEjXJaI9FxSRh2/UGK3z5Nsc8NPV3Htu5LvZwCAY
mM7PqW5S0+YnHRLMo4d0AW05hisNkPj1j/2fv3IhyHT0XAmxLd5ZvbPu5GBZ1xBGzWgNtDHS+RvH
7fhRXbAknubsPXEMfL0az9IcVKs5na82JSSzCfJ41tWtwERQ8lbD7oESQl5hxu+F95NckKhxljDA
JN0oUYq1zQrj4TGYiyj+rRng+7Hi17lZOwKGw4iZpd4JmZCExd6MUGRd6Sox2z5X9JM9N31O2Eag
pNmK9MkeFKBk9gd4HIvJJn4BA884qFh+GXBkbDLY12JNK+avxdi5PAfmLl8vQbn1MQ6qoDGzFc0R
luCDiWrxjrGi6gmVj9hbIkfnpYt9oPDYu+miTUCQne76VtWmMWbTtkW5sUUdrOaMJmuBKvzOkbWU
rbsJVOYISkfQiMjxtYlHarnUyfC11Rp4w2d9MQCkihHxltvSQBy6pIOhJ2GDBUE5QZ5OcLTVuNrq
muS5B4Nppw6S6ZDU38wF8B45W6mbGhUG/8FbXNaad2RHs+sG1POBn4YIWJSwZezwWCph0V66fVV6
M08MHDw2tbwyXEiU95VSGRC2frlMNATCkviVwt0FEYaClHOFPylDRHwLymMjV/BqENiPsprf3uX6
fEo7LTlixJQJ/QoeiIO9uCrNuyjEKsoD091cxJqlVyrru73ojqmtPQ57F/9VGwgBxNDf+ASqyghR
5qJomW3HUGngciChUpFWdGL32rW7b0GshKZTLzpHQVVgDLQ808BAAi8k1B1WmDt7yhhzeWe2FNOz
7AxWswW+5hohx9oahJlMVe0azZJ3nmJB8dMztbKvPTU177AdtXzSYthNS29jukuGTGDez0kNnAoM
GnTvFGmqILZvCxPaH/HNFRYjbDjGYzD7tx9hnLFnBukiCV9woG6OVDMibU9BNswaQa5Is5NuELAh
tfw7xdBoi3mcifscs1+Q3Hc5FcgC+RiPX58uq8G0fS6I+D1GZo8pp9nnil8fVsuRnIFAc7sWWZC9
pVFVwL3tJ6OG9Ik44d0QMw3amGdRDnkCDvLCVnz24AwRE9N0kvNiJe5sp8kHoJWpCGtpkOgw0LkB
dEMwG/0sP5ISul30RhW5JJYjeZ53Da3OPp1vFYGvzdeUm6cOGOhR7zMei4FIFFNpj8Ln9xInt4VV
RUD+cfp+ChsFFE1RC8/TysnN3aZtdFZYV6VT40TT9OA8NunSSO3njsIPQ5nCzypdSTr4wYQ69VR+
hZ2/zNkMA+OFkwiyZkmc87xjiba4HDEVt/XFAYsBWV14QYqK6sGrDJo88uSp1R2vOMvYDsXG+dF9
Pgj5SfF5ktPH1aWKPKu3fkgNHhoCqdcyX9ZAOXmLP+jwxttlGGgjbzCh2w/k48TBb72ot2cEOLOw
AsWvZ89aL7NqeMDqjRz11zchvCXbZBXgOKGTvvph3rYZi4mr59GCc7Swx0RtJ3QgFgUOxMXC5P4F
Z1W87WT2Bby5GzRxNLBOVJYkbeVhQ7eoBvbdMIoBYockuVkBnK1ifInwBxbGZfVw0Sxe7BOntd8B
u9vFX5SUpIjmi8idD4P7tXb52Zpj0gCndDJWo/+C3HftfQNJLwNbB25xN5irs/A7GtoVQWK3HpcR
JaAI9iqeObnY5dPq8ziwIKTm5TfxWQfG0hQgBIwWHkKbV997uz821ECKn6ynKIRJ8M4oAv8ot7U3
5oJYvfZcoiyp0k20wx2Skq/J6fwF/OPy1B1eM6Sf94Dj++3tf7z7xsoDVFo1ukzRb4PGgLVe2MEB
/xvv0ljrVdr5GTPaHBSudvQfyu+0YIZTId1jgAXyjvu5Nb8PfufUomN9Ek/3q7j7ElcszSCq5eut
pirbH8wKI9sBlXZav48aB3plAkpnGVWGr3R1B5COCpasrVYi7wUXNOp1fsJbJ9j5nlh2LFZuyeIi
CP3k2JBxit38KPvMEKeQbIx2uLwYbOsnuRl45UIPUNwn6lJRHIX742zByiZU+7VuZJyxIDd0Ghfa
xjnDZ+P42ORVXN+EHx+0+CAjoIXThN3jnIueDheP/WPmK3KYxwkv6ZtpkT0E/JNCc1FX+sK13cXb
B7d3zYe+ypCJK3BUuZcVjRCYO8cNBZxjr9MdKBagPNokSBeKJh7Lf46BH07njUBc58RKK7KWCUck
+9hg0enTVthseeSMz8yfxhSpMngc4jnBzLg9HjBi/4x904XspJWXItZE1ljhNkCQ4ENos62vlG8O
WQ1BKa0d0qYNjb/4diW+uZuGmh72b0rKc0AtMJ97e72UkRA83eDliykQPHi7zS66CUkvsItDOQQr
ZyVHjnVabXdokxHpSyNoax7rkxVuC676bdSzvJKEIWz9IVgxRrSEf8pmF6+vhXRneNs1OI1zbSSB
Rf7LgF6KPam/FsW/xUJAuHmg9BUJVLFrmG455P1PMhpF1kMqm1+Uc26zAlnOUCCgHAexBwo61iOe
ESsJFOkK2T1OHGvEzvAbx8MVOZCbnss7jb7smZLhvuISqTFNw7qOPusOoiERA/+Cs54vaejxUF5E
0KIN2HCTq1x7qx1X591q5Cuh7xIXFmyPsA1Lvqg4TBepNGOv5GGXDOZmfGMyNcpMJizd1wqsslID
I2haO5YmurZhL4xezS+rbq7bVMQROEPmnmeq4AMXNvQs7H0mn368EN8Tin5jFX1NH6Y16cWyf71y
/s45P7c5fc1Zcj8Rkg2nC9BNc5Z7AtMQbPBBgAv9n5gEgAKyw4TjqHCo3/K9jR5dzVj1IB8T9wGc
eroYJpGKUJQdr15+ZYpChjgXNa9gd70DALDVijjN7x4B1ZVsSKJSEiEAEGwrVQfKPHzJsUGvNQbO
moBIOk51JkhDCRAyZwihC+nln9CPVWFdComPjE6W9agtEwiuT3XUTKTZpBeuQm2zIE0Cn92NakuX
PAzB0PV05OLL4LIt9ZRQblywHTG/LMjN9L1bVlDKYw8gHH4gNEsREIQWokRHug/3QEH0OmQLrQKc
lFBIw3gP5yceLHZi4+5AbA1MCN+ASLxmwDjGDMfw5BlQN0JrBDwcxEbuZIVzEC/9X99vQMSzvT+y
jvWbKhcpbGfW/aX2oD/3sa5GSaOHHWxAzQo+ujaJKlwRZGuxY1fIf3hxHYvfwh41wdF0c77KMWTi
VyFuXPY2Y704TvTm5VBgmV4ZkrhryRgLWALlPTWlRv1iyYN694RpJWjpg7XpPxl6eXjMR3ohRsku
kAhRXUzMxOtcEhlKhwA8k4qwsvC9ywHmYNbqyzCk7Z9y7R4VQ0LJlXz9do1T/vkaiIDf0fpdKJDt
Jj+DQLE8niGPRwnJOyEgSpIM2i9Mq7Fcs6i3fiLG70B00oTk4s235e3MpdZc1V+0CIGkeqS24Xfk
wQRvNQMJF9zhjFqbg+8+WKyi3J4gmVCVqFXv8r1IGJ4IRkYSWUQPHHRbxJRh89p6OkRBqCW6mYfO
NjV477hHYXIMQJLSKQJ6+pWEzCNTPzJ8F6Cnqhb3chXQnDUNGv8dQcphgS1Txzb6VG6SsfbyWdPh
9paw4egI5S0YFtCvThvkq5MEl7oxv2zGTJnrnv2sZiLaU08+69P0oyKPMmq8tKLsNfUOdKQQzlmb
0D7frx4kyJl0Srd4yqWzTRd1P7Swd6BIqPBlzV3cBqoa2M1ADSF9NqEcggs3YVpm34hmbnvliNxp
TYDExTGoi8l9CltLwsm44kOuQyx3Vl99QFarOEFaFuC3HiGpkCjQhND+uODXWhY1QabvJnpcygQJ
u+rdSade9e+0uK8CHPl6sz6ko+gP2EzCA6ET0wSaMf15IxdELZnH04BFUPmQqbeHV+UOYMJiLOEn
MMX0VBI0TcRXiD13dd/gIGEtnvs+gjE3LjAkTAVoBDck1HGCTfNxIg/I7AZWA4Hua7QieCI2a9ng
ohNll0hyLammK4E5W8navxw/ZrK21eTtyRHrhg4g2GbUfHpWazNuF9oiEk+mg9/HMiKobLf4IT2A
VWRyQmcEjOC7oPrV9sWqUfnB8TiwuteNcf7ZDGLXzuNAenhaX5i2TubwG4JMyWyn8sukkyYEDoOh
runQIrYzpy0rE8I8NyAAhjIcJqqwJdcBJJP6spr4mM1KhxBHj7mdlQI8d6QkYVJ/ehLVqosuKROa
1h+mgaKqMPsc4XQDK9nlqrF70B32ZCH3jjaCa91BePRLuNYmAASPpYgW0BGr1Wb7P4EsLYOoCkIB
TJ75IdfewJiyGQu1QgzV6GiXqDY12EWAAH+gRfQWNN1gNOYj41l4NAAX0IToJwykTlX61vVO+pOg
wI1iIs1LaqLGyENW8FgPUvaXgHZvd0TyAjPebOZs5Jngk3M2sbwG0sMsXKqYa9arN8g4cxh0x8do
IBvKOwzx2tnyME2ppGAmRWKG3vlAcQAmV9vjc3X/vXgHEzWmF9qoEN701HdEvmHUM0VyWVZPn1YE
Te/xPoR/iNANMap+It35AmshLq7C7kLIuZFtVUYJMhjC9pRRsNyG9m/fOFSX4klfdmolhOsEUbf+
lzQzNVhJKgSOB7Bn6jUroVjB+EtKuwNBBVIisSeuNoIEaPjw63U63uDYjs1r5j0eGa6tCJAl266+
CnqnVCGzq4QXMp+lhqG2f6VqwEdaerBv6RQT32irhqt+Y3jj8MqtBF03a44siUw364H94k+Tgo5X
jbl0/GBUokLj9NA9zb9Qn5pa0LjDOZ0quG3W3dXjrRBQzUi2IiauWLpj3a8T+ZYUfAVOgqA2hM+d
sGEIRVPB/uWYnwtSR0j+Ax3OQfLV/7QqTgKeZkuA14h2LBqRfmNrdeuYr4ZwJx/OyulkU1KfZU5O
cYs9elF/e57DCCv8WCdM++fcaDTF5c3ypzNi99N7xMEQI8S6Aj+jvuhQYzh8odANPiHqDPRnyEsv
UZ2rnMunmY9XeG8CyF79uffQ9uj/vLQ8hqTx/1WX/jR8gbA2tSZkRJX8qoyLMYGBw05CY//q3tkq
q1dwuHtSeTs9RJosInOEQQcwkHOVILzEcJhn4AlACzDxytYr2/KA1ZIFehaCAaTQmrK82GVDlAbm
BH+VuybXKu4zU7C8kq6LzU35KqQ4oiVFCiSSo1Sd4ZRBZGpDMy3+KjwVnYLOyGmd8Y/8SyLjVKN4
rQpzqDC4PQ2Mo2DUE/SSQYc1dumNLsRuSivv9Ie2icbe+U99CElm9s37dYR47OtZBa4OZ1DhBtfE
8qPhOMiqMrQSt5tu15tjGgHX7tnBfL3Vphurlo0HuMx5szSikMUNh9NBPnaUbc4FOFByWXov3/qS
W8299H2hNBiiA15PeD2HkJ25CK2FwxKzLh7qI2JScDlPCBPK0Nx0TWfHHc4IV4WmHirNpzRU90qn
sgA7uzaWZKuS7jfBgjaPUBXGP9kbfTf4qa5BlCuk6vsxXDwBSOrXo4P5GMtiOd7gHcC2m8IV6+h2
4KK65yx51zpwl9kFtq4wy6y0Zz5TXvmts835azllHsj8npo8UELKD4SNt8O4A0l69T9IR6rIJ8VH
IWC/AdWruZBxz2SIWkfh8u4E6eHyXlUVxHfghLmCTM+Ivn8jNsXOtR6ptAour4psp3xdjd+BOWsM
auONTknshLaFVMRncMocxOMMYi52QjPBFOHBG4p33mDCHkTyvhAeUd8b959l3Kk0TRCegz0bqsFq
NeY6BzLDjBxlPcZicIUp5jW3DxSjRSXNm/Hu/TkqKCI/aRJYQvHYid00KB/wZwbI/9ez2XBnr+px
Z7w/x0m2oSA+Q5sCniIWTaLL7uEYmakldEQoneiRpuY+7visqUYRImexlvdw7XmPHIkVRB+mjZVE
4qUUocKIjoI19BPt542S7aAwSqBtmhCjpQ2pw15olGeFCFsa7jfrrnGGbpyTdw+qy9Bv4iAOmJj7
ryhcxrA+nXNUv0wT9OdR4Qd+p3QwhNHA829+8LVATfoECgGc53rms76b5L6tTyh5DuXZrH5euFHm
XAd+kbYi2wVbpJQEPHrUh87wplx96ArFydKVkyVqHyBTiFUIfpHQlRpEjxY8w+kd/k27sDJbOgse
ZwO1LmaAsGY8DLSPZMee1NyQAZBteWZ13kXNLCyAP65ShPjX7BO1U3AvsKcnSUI2IqZdv26Y3FMM
c7AX0SDk0CNhYcA4/HedUjCB/+HzamLYBphpgOxghKPI+39S87vdoVcUUWqJqdJCrYeHS4EUyeWX
Kb2+RbjDWAaTQYqELZC77Vvx8Be0xZITOV3QJySHrSqaBhPsXw6hfzfI3WLC+wRwAm5db0nN6vGY
8vqHYBBMbMF3rtlG3XocnSDz2vNklJX2lHwbiZokJYBdcFmkCl7KXswFHX/A53oAFYSHyvLPJO++
mghc1O+g/V4qF0rTNLdoaF+V/GGQwe10wuIK0PieOyEE2RfPdV8Q+cI+F2++1Z6HMfjiz92rofzs
pUbmUb7PAvKlrEKiXGkNjuIMmaWqt4b9iWMe+EleIHfSS9Dm2N3Mz6lj/2rXZ0SAjrJ8Jp8hNmUC
Bj+YYNLwKjp+3Kzu4p5zY45O+MVu1VBk8fp8pEnUwT9d03hQJFsCcRY8OSW+kBscdc4PkRFvTMfF
a+zMXV1B9bVyCygiGo1drzihfHywca8qkqt3/+QYl8IGvt9BOpbA6wlwsmX9rTMf72vncYJTstNA
qUt69kd7EI//3wysntejeztrMNgDkqG46GlzieD62f3UtG3oaVXrorfPlzZjAw4mB+lUdmVhuDCr
PbQUKi60xz+xYVPBFbHqdx+ZLHZrJ9U/idDAPrcInyPA335vLvPCANdug1PjPixqeF4H24FRojIe
s+ScCJ+lLhfqKVG+Q5rnEpiXmCwxNWZyL6IlfYQBox41GFtxs9I7233yab3Cd4LP4UqySTaLSdDd
a9tmccAvVKcnFKLJ9kTk0nrDxxxfXVJz13/nhcsQQ7po1vXbA2gzbcghnfhviC+n7i/GTp/IyJ88
k34tMGojWlroegp5QCnA/I/slm264uFwRRhda3NewdNg5a4VwDfO/AV7dMuOs5KB/bmFG6HnUnUk
dhj1aoimBAFelsLDY6rvfQce7lG3EMz+eqDuygrMQPtSBs2HpysiNQcu6VDk6bqt7VDeoDMqK63Z
aMQ3IfbH5Jg00AVCXU3wsb0v2JYDDKvv7OFAyZZRB+101EeSe7LMB/UqKV7n2HZaBKy5bY0uWyv7
x1vkIv0Q30/xE+KiWljH7Nw5LBpHw0ffvx5PS86lQBmguntosWZSdKkbx73gptfYSHfmP5rwU41x
LvqzCtLys8U0rahzLTyhoocGo0esK1pbFc+ucP3ZiARgDY/KI6ACzjIjcHoeibD05zPxLah5wCmQ
sZL6nw0XS6BjWKAFkwTj+1vAXZScDfHFODwPyKyZDUDZixkFufBLIkpDFN9f5pqEKm3WOmbckU0z
rx1x8pJGFzHWWGK1NIpYkaCbcTLhKI/pjMmd1QZWGk1RINMtxD2evRxEbvfCoyFBelX2VaH1IqHI
hitTSti2w6+5A7SLgNiPVgnNvUkGafTGOotTe+JMJGSFK+h75X6K8g2bUlSqno9aiAowUhH8CHgc
JmofzLyf2OZBmyMjfBcnlRWXpr5VJvg9nwHKMU+PWmQFUJYDzSjHO2y3+3ZyhzEtPEJVaXAuTW2q
Gglg0SFe6xZ1oV15k6/d94rpnSyK2aAvTMI9hny7OSiA+a8ZTRzU7zBvfsV+9gV2uGfgZdl52h/S
/nUGrHbC8QqAbStsM47D0CAgdhlT9RefUFFwsjE0js6xWBjAcXc8Cfaqg7CeM+OZ6TvnyNBHAFIq
kOfphyT2EIkBMDDzBYUUpGm2OpuFm/4OggFyhfGRx6WNrpjpX0rmDmN+8/BpWJrGk84/pWFf6n76
KcVlPtsUjyvcwhB7FTYNHMi0Td8mNw4gTm8YNB7ibjqDZIFJCkr7Ch9mIroqwM5IDK57R2B0Z8Fo
1fuNWEm1QplyLzrXFF3F4r5LUX5Posg3fdTTa6q+oK/EtAaS6XH5n3FSZ77ru4tt7NZnAVU47YSq
p0V+gS5p1aMXJMNjScbbcXoChHTYMxrp6YHWcCSH8cwktwO6qy2Xy8HiA7p3ACrhcez+RbLh9YVg
2v0B9dDyg7t6my3Xt+1aAWvYIpKNSutoO63vfZ1iyPnc7X/cf8r3wLjFmBb0FgfoY9OVugg6Ribp
ud7jrYHdlLfn4kbQF9IWcVsS/GKcyS3NheDdamHnmyZrkhcBCaGeWF1dTpbnHKVCKl5HDAc7+EIL
BcDxiWSPOkujQ00sUW50UxO3n70LFaEoL9pGWadGepS+3npop70hZXFMNFDBxfeFNHeLGIsjgc11
fuN5QV8VIz3lNbUwhJKh8iI22hPx6OEfGjQ+ny6hj8dJi9l6fQlogodoiGhiZZi7ibk0Dxxk+zGg
y8ZXmqVl9Unn88XBdAy8tzNRrvNtAyaz407k+aY2eltT8Bdg6Kt+e7S7PToVOiMqiIkAE/GwbpJ4
/sdjzussOt/hz09hpQvri1opAKFJt8gUNByBD9vbcrEnsWSyuJ7zTEYTdg4wZ2plqTLNDdqX1QPX
ZjZa0dS+5sRNbNWNiLoCW4sWQ0ZwafzV7ZuZ7KPEPbIHNPu8EDF4TIoAo070TXIlh3JSNgpS/Pto
4bM8A9FliUW4Z/yFi7vWggIILVlep5dE4UIvhQCa7+buUJPfksNpM4x4PkvwhGG21OZQMH4ewCr1
1//hvw/c322Q9QDniSgGVEg9j2DZc4q+b5Yieii5E4frmFKjFovsnJ8Ynb3pqSxx1lhyT+7MyUxS
NfWUv9v7MOJALf3L/tflR1T2de6AYl2Ltvr14a4ZhNXIP7uvYK8S304NosWXEHD3zaFjtXXn1z7Z
XnZHpMiQAZty5IzyCuVwOu6oNynvR8Ee7+reh1PzcRuNZL/yHqv4fOT3MGgIrGPtokpDtAtT9JEz
l7F7azzSyaOyizy50h+xShBNDyuFXoAlZ0LgyoLegtLKOI7V6hphPTtAOkdJ4RVmE8I+tPqy3cjm
0k+vojoFyItTT2Zo+uaHkBYUME5jX99JdzKzuYcyJ6y2d5yYaWlfWh0EMk9V16xOKxoXzIJj1KzF
d3jxhbG5uR3SIXrW57wAxFMDEecWGmpwAjfCeUqPRH3CF9K57fqCxurW6cqmdbmte5moMMuKvfdT
1YfSMuasNGph4/wpc1BTm/ZGey8Bd/GXiMyFO3/KunAGqLUMkXzaXle2C7aASyxYaNByWu9+HbCN
lN6fIGHfOnrbuBdl6F7+y1YJSmpozfXs0iOH4YjlYRaDMpWibMKrenCgv2+MJAAqWNoeXUffbs7q
VbVKQDyBBPsGruboJLSo/3EvV+47l5o75SDa9jcAw8IhTpQtif3nic4/qC5us5j1g4T4yqoq+3IQ
My2iUcf1OJ4TKBT2bTb+76RTczo7RyuDKMGICmymoo08u7rzvvu6S0mYhnfpLvuFCAdSt6A4jg9z
FLF7/YW2goYyIr+Y9gm3Hdv0mbVhuFRyHeOfwQS4c5TGZvt6n2vck3Espxz12frHVezOeFmjPAHU
03yg96nfUXQYdt26mfzYUmwFfaez20DqcqtBQyAIaSyVxIx50UlooLGDrulCrEHICT8IT1oxSR61
cRz38jTme+zRRzS2cFcJcQ/No6j7HHjwzPRUIa0dyyWF7K2TcY5C5gIHl64J2KlfZDg8GOop5zTO
TLmHGotajsXiHDrOvrbKvP66L3PyFalpR6OIvMcZ2u8mILNJZ1Ia9x9I0VewEY9ZNc2OIJN8yBjO
hid8XtFInL5W1QZxBxeybd1b/gygbld+A+/t/BR0jvLyZxC8Y6mAH+2p+QYeJdzTX1C5+rGsXzCu
7ITwOksc9autljy4VKC95Z4bskOrVhTXMT90Q2yI19dcqdh4ZtbhqJTJa2eyfQh3501WkrG/n0kQ
N7tv3s89/Mhyj+FiTGChmIlWa+it2pUHijgrJYr9IHr2uewRhDdAaCmYq6B1laXh0PrER4BltMX8
nZXCegagNRGJEjH7RCSH0rXh6SB/vvGQgTH5hrw7/ArTzE60PFvW0LxEK4qVcmaXCwriffcZzD6j
ynOT4r3aU2bMt/twjA/5oE2l8izLrPvmMAFHvIwV+jRgkl9i+MeQTEh8jrfbAzPgBNbdlb12Ntld
8tbet7/UpT97owwYY2ZeprTGQuyQcW/nZdYSQW3I20ef3IuhBhYIWQv6BmP3SVOi5iGoWxzRdfO4
BEjtBIn0RJO6d9KaPtERkTSGIV08x7lr0dSetT5RC7nw4E8j0Rm1W0asp9kDE7/7e6/MusrzlFLe
FxjV8Qpqr5iPQKXSqfYm2MfiSrAJoEl7wa2J3BODJ28hr1VGBxbtMmM54UY/HMKUNNfYIJMmWPQL
bnFu1pTbI7NIQ9R9sWRl7WI0y/ljTTihvMQdD32tGfYkZQDoF9C2rKEL8AuOptgBhhmZ+UOB9Nk/
/zyHnpdxaoumsXN7P9ADQPqR44+JaYfF9KF8uZx4gWjVzmqGFtZiaZiDcFa/6LG4Xb1zd2I4EagN
GzrmGbhUE6UQ6G3kIduWLGyI+upso2lte7ze43RE6WQBGxRshRwwow9kqHNRvLYDPI5sJxkC2gBA
UU0UyJA/oZlX8SmOKUj1Sqlx+ppU4bquKnSCPzfV577cuvxOJQRsKMW98BxAeVjAVKz0m0Oj2aRz
LeuXrYY4tzwF4QIg6adezfvnmCk5wmDoGtdSfWHzUM7diubMGL9/vdLE2QhehKJghWOxT1lAcTbm
IwKQlL7YkmTyt+UlSxN7vxHTlvtOQujp6jx7Gy3E8B/T1n/78FKAeSzbeVdyJdYSQ7tnWaR/KIvN
vXKMqP389bibvwAajQMmzD8Hv2t1M+pwKc9/sFAifizvs/JfnO8cGfAVkTvJerYVb+Mt99ZG+pbe
TmLU0SYI+fOEjq6eGZMiSo5PpNOyKsl8PX4XIpYzAsRidACmlNYlJfDvmrRFobw2NBkc+62nyI/b
ifQbTOTKZxGYdyo2yBRlINfc9tAyLyjbr7cmYLUlUyVh/v6kpQ0LOXSZAjZvSUKcDALQ4S2s64t0
sLRZchYWTIppc8AZdc2fEqkMeqCb+vssOl8IEk758BzBfZkIQHAql+6nR60TExr7+77xpPLjsJKH
egAaCRr9XJOwOXi9/rV0YS1oF5fWARx/y9SvQRtx/ODGTS7RlB50pHMxroZn0yvT63xVeoLZh7wB
TsaZ5zp39g3tEel+mCKPDGIQJq9AoiIEeGXyIisOFQWYpg3a3qZMuplqnacw3ZliyUS4M1r721YO
KSnbpKZwQ9KjT+jEmVtz2pSlXWqc2qIkqxttiiz8ojcyZ4wANPK3EwMoszWERYNOzkZ4mwnEC5hp
aQtoXif1rYsAehiVwUFQboXCmOvl3Q/lMlFanOrHID3aRg/I6yMpMxJLDfsasuBQj2Ese+2MpmwE
AT/UsquMHLlWUdpx5iJPexKLaqtCcYOeo7tsAraNagWcaZN4tUbWV61kifl8xVT7/7FBfq3lL/iz
1z3gZTjoyW/jKlK1RPDlEWJSlo2VZgQZUM1jCzSnxc6DCwuCaxZHM0sbHzRqPp8T4h0BCTF6lmWb
sE78zlQrNyfN94Cc+zkztNpTrwmIRjIPhb/wWf5XdV8DPFbNqVTfeoT7RAMb1EWNNvT13zlgYejy
2/jDHjenj2QHkGnIPyP9WfdT6Qh8nh0+B3p2uuIF96SgpqmNbSDjmsCpPm/AYgr/D3yNwKo4S5ae
EIpvQBN9aeqD1gtUcKlnu1mdZ3qDi5AFqhUUqfmJ/WEzYXm4JZfM2TZo31pKwCc3Qj+Mkg2VC9/D
mEu2RpLoG50RF8G0ZXzdX0lx/09Hq8rvXY4sCKz8Jp2AQ1r3+GY8+eUTmNc4Y4IqfwJ+omKU6WdA
ecqJGGigtjg7cRgyl122GPfWpUQtJ1Lfxkvo0ltIGyqJlhD8r3sXgFXFKA7KJnyidnmiZPhrx2WH
8voH3tQQ6GGpLtKk8Eob/076C1m1hTtGZneMqFYps97Nw2A1UTNOr/pZdiM45ywL+tB7btEDSV6G
nthPOuJCjntiHhUINdh8m5vPv+Tnz8kckI9r2IvEvOCZWIRyWXweU7qwVydL33xog3Brba54R7JY
Sni/jyplsz/BZ0f/NNi4CmcTDVz5rTTi4Vb17d5TbfiJdujBGAVaXFa1TPIlq25e9EvWQPVjsQy6
6MwbXzOJsYBmy0iIUgDyJ1DKF+HRvbOc4BW3LEv++HefUIrX4LDTFK7rrc7NoFIC/GDTkRtksd+1
nMo9fOYq2aeyFh3ytQJmaqaYjSCR3u4yoXVVT3PlkyAmtEsii+/itx0xKsllPQOVIIdUnruNfblo
NQ/vzKQC+FrKcxor7zAXK1H/ZVeedlKLkqDl9IsaPyc+0jbxL4d4tcuexJJq1nIxy3uiyyz5Tiap
ky7pR73/DzXCA2FOxbkCygo8b3RpZ2tX3+9sXfnZq+DfmSM6YOGPziS5zUMppyZc9osdH9P2GqIS
n+EYF63bT/igzwAgTjiacJHn4+fv/aAi7bEU8GUfqY0406FMxtZWjCGQCsbBG2l7SL8swkJkTjuu
9xfurHv+Nn6Q3GQxxReO/qDesqgNCYjsWyWMhug9Ihq2djH+l66hnACetcOZqWj1Crh1gGtYdw9H
GOG/LO2JOpbqIH+h73O0uiWVDDDc+g9yAmhQh8ufcZgVdZhFW0gfJafJ0wPNRvoFgTr2O9HA2tMD
An2BUwMGZxgZJTq/XTOxcOksffv2OVIgRvA881IH6Y+Lqgv9mLOKA21enMK9Di/JR9PuBpRmSWGu
q2ry8dUkXrTfurqLFh6eFJhf8Cp8A6SklAEp15sgcfyOdqFTkWpeN0zXKg5350IioJEvZFvPrWUi
8aNlfZ0ATJS8NX0pSEr0f+c6W608sxJwH2m1ZmXzVYipXzWptC0kuZdOzot5lvK6aqZHWrX5acQi
6+isPsUJzR4MQiV6Fx42/1Skro6JOi1gvIDCAQSX0NIm7FVdJ51Oqj1XmgC06BFmqLOuIcvC/Dj2
62iJW0rT+KeIzSrM6DhUKPZa3HaqIv6jhwdcIP8FLG1snz7B1cnMW3rv+V2y2ZJCem3oMho9fM0s
aWbNFzwdlafIdn+Ta8SwIXSKXPqwfhk5E36Q+ZjR7PDTLEpR//nMYql7moV74vGXbzE+dbcmN1JR
3K9a0oFoqbnIKpZkERtEJKiDVrKDG+PoGA27aujYJMwbizPpH8jN6nc4FkgVz863p5ZnSkQoHsMS
z77OpKSy2FnKJgPtktyGfH0jk2uoIZzSLMEgOmpiASMu1D6TurIdz1NYD5IbTKeZiikBTqzisy/H
X+DrvB+8eBK8ONJ9Zn+A+J63NafOLVtd/Kmj7Kgo4ERGYDB7T/sAh8ut4+4IUDQ152HT8tsiKWMQ
mEvrO/wEMGXF2GRWgZL+Lqr8Iw643R9EjeY6L4n2bv+GmsOFPfmdHad5uClpIP43nHbP8L5hU0sq
CWjC8eez+tzLeB3PWal4PKhvsLIPYphmk93NNlDLQfv9ICqzYfq3GJ161rbUHSBfWAasdMAYOdVy
x9bqNXQgXmKYCUazq1r9QfNuzLqOX+HTkKVjiYVxnpFuGliIC+orO5puoW7joTJa6raw3AkliLWZ
tO8CRMp4ZurGB3Xwafz3lD5qN8GzHTyIHcLROI7EsUr1kpPoiOL+T7tqsGz2m0offALwbfBnPw+r
2//UbPfghtAwtIPBdSlPQavD0L8rhttJqceEkIZUHMwLUjt1vs4T5fRsbDzPEVyU4wnmpp6L0Vde
5ueNXEvbE4YKPKBmzCR3O9AEjB9eWfef4qZa7pdQ9sMUUIVQTGw2dYw0JCrotI8B+Y5jJMwUcpDU
u8pXIRxYvCi96z63WTHksfDxhCI/XTm6blZvD0wjd7Va5Jj6OLrtkj8/gZfuLy4tlisP/104etkI
5lxPDruwX1sX6Vbxj99pHFMLNB9MZMs8MPD5dSGQ8g/e2zGgAbXiL8zAZ8FZxjklrOfzr5Sn+PuS
DtPAhCRKxsaMrwTcFSr3UvJZ3yU4dG7MzCvZczboz7qvtINFO2pO4CvSdOK7BmSfLMdq6oFABVYc
xQF/MrOzKljds7dFHH7WWk433niTTazI/UOuOky6EuowkaEsV2Fo+kmL136wX5SNP4Y9bLvXP5jE
RT1J7XznW82rkUg80bE7nvHRXWmz8XPwSd13R5RoE9uGVwyLU2y9897N8luKSsALZYziUU+eCyGW
gxfzN9X/Ssm/E+Uh7asYsd+bFxp7C0njlIbDnh8H0Ma7MjtJnt3nLGQ/wv6SJU/vHP6unwrpNFpQ
k4ufsABvvDdciR2zVKwhonrAQwYeHS8eYHgJVigunc/Otb9fVHPYZ2gCUXBQhTfMVv75Ab5opEnu
ul6maIo0SFuzqikPohhN25PjFpta5rVHEFqFEr6XJwvKon1336Es9kCnjo4srLdfpJBIxIz+XVGS
ZY35yfZzLrQj63e1LUF8FOeAuCWx5uXOBmElnYn9IYOiLB9tqjWwVyUglSJURPL07MvsWtNbrU9W
AwDGp4tV2KiHyzxXqZLp+M3PAiybgH+sQ4YRwU3N5lhV5XP9ot05bmIwUU40Rp97N4ARSkOZceZg
UQlBJK4VBFKqUze4GSfcUOOllAohIzCPGs3vyJYIe157tqFMXzC0x35sIe/Mv9kYfwUEGDkfWUsn
MVYO8iOzKkyBSlYMUgjLJMPVKGKCboUfcTwyiEJQaDvYOn3uurFYFzoSma/ZbTntQBqx0LMrhyP7
xEkWddca5/6xcemAkkANrRb1pS9EQnR9AO+gfC//7ETtBk18lQv8pnq7Pn8QKSTCRpS9Wo4JBwiA
yvCnIrh5Qp1ODydCg3rbr0+9CbIKM3dopK+XEHUXzu/6R60lay53c+CrHrim935KvH5N2KbdgNuh
qZgW2x5chyeYG38PrTa8oLboXfaUYBqag3pPtTIKeK/x4pbgeDgBR6ZQy+gTp30tg/3CgYKQXxHB
a2mqEw99Tu0WomrgXm+/NjMi2xKD2gvZa2o2wQU8AFim+emfFAKreNq6D1hhkiUsSnO2XNMtOhuC
4UIhA+ARB6A6RQGAQEeZbQ98kKyf3pnRm5/cVpstJ1S32395BLupz17ORtD4VHmSwtwlRIOEp+yV
u2ukAW+83QHfpdKYWWzQyBt6ULRjBmzBF3SBW4rIBwVvSL/yrxkpAzGzVYEMfVutwf9X/3atH7e1
H3GA9F5M9MK2XpIhQO99Fae6z8sDGoy6TE2z/QvSRdtVPRvGVPwSGRFehYwmlIncqgwdvOeapSn0
VB1FOA/Tpb1e6c5+uOkIn5u57awUtLCb2IPjq+rIdQCE6ADetZ+DX2vMJZvTdrRRmJQ7HU+PF9X9
ADSvTxakLPCGcTkCami7NzBY2GtyKYTDEoOlp1mH0+N+iOnOgODwC6yRUUKZYCrLQuazZkNND1Lw
d4zJJkBY6taa1ymkJuzbORBTdkhS/ZOdMX1yKocrs1pidcukcdOY9JAg57VJzD6Le0jj+i+TTocW
AkJr/gqUEqVl+6p0WCk/5x7XmP/yXn2Tvj7+S6+PbmH7vE9O6UibR2jYneLiw2GijfNkQccZrgJY
lHXQynp9tbSMHhY1pVFHNxtkth4Ibfx5+ujZyN+q/OsP9WliW28tfk87FqjvjCwHD1cUpQ8MGlqF
jeQ4Ewy+vX2bR7oa2Ihtd7LaJlX30YxSjpXsP+t07hDi67wR5VAISU2H7XRxgRkoCTt3BXZ7aYnd
8/rlPGZg8qncdG/XF7wY6LbaqRMsBZ3fysfqxmPNT35pbGpCcaAPlY20Z9VATJJs/qW1FN7zgmEO
lklEwM3VtSz8E8zKIu9neF1+eWOyehFMOJaG8i+o64g4nlkjC/AVndvzGVC9SqZH69yahiM3+D/x
7LPeLTxOWaHb6liPwqyXYlk+N6VxbJHNA1TSrAnIowq8dRUnvDfI9ihAPEGQLS47TrKFyTgZrJXW
4ACEp/frSCYcYf+qnmRAJDrnqFVagAmT8RCHwOX/+Y3DVu9raDpQAMNqgW73EPOZQjQCJGNjsT5h
2RTTl6gF/vxdCd8/2ya1oePfYipmf6e7iPyehP5/rSuMLnVqbdapI1JGgnlGBWMLlaiLUmSbTDbw
SBNsuaOpZlb0n7vQuDeoQ7Vpn66tjI0frCIFOIWdUZdrEntBTXrW7n4vBp+kssLpNUAsKfD9ccS7
nDd47d4ch5QhTrEbt/e91t96D26U4IehZqI/9dHCs3+4EZLAUlerSKnz57aHlaacGJuLk2e29KvM
3FXLLSJT/NgJ+hRbxwvdqAdkaHuQItvRu9mJM264xlhw+5gFrCK6F3LrhuMw/9lP4fmzZccG9nSF
kxdFQPOqRcV2HEoa/cax2l3y9V7GvCGSmMWySeR6kvUuFGT98VKyMNRvDWDdzPgz+z5fvz9WYnhw
MJY0T/Rec9lMbnuPFWv4djHDHavwWTjFPbQEoImYid3PQ3OcQPwU/HcWO2jxCJec7zm8yXjk2DGO
rsw2NHU5y0U+Xrgg4PWd6f66xghKnKGbCQCh0JJo3RPgJ9LXJ+V5COmk/L2hiF6oKWfLh46KEeps
nQWo93vx+21wymJBtGZVUlqkSN3PE+4OSzngVqh6HU1COI8+mRTlont7nngSW4ZA4dPuFJICRMg3
suBguJCcKVA4GXIPD5PrD23XFblIzy4iIwd4zrNM0mvCjENEm505nMUegmV/nekVj1J55LGEXEFe
H/1VszZ5w9foCVrV2xxNCcgFD+ya72DbLMROonKfc16czr0NlKcT6RvM5BHBYUYTIv2X9rmgYnx4
MS5RgSH7YvhSTirrrIOO4DIL9rPVP6EHj8oFH5Db482GehYB8R6Xbq9swArIU2dDQ3JVYgk1O4UW
s9iCtNByEH0Nr7Wx4Wq3kUN3VacvZQjDipyFMucoqpBE7bnAOTKNfp66SCutZG82g1z7MfTZ5GGl
qnzl1pbiqj4GEhJJDBdWHNg+MYw3gpOW+Oj6BOymL2A2fIiLoRmwp4OpWR4XxuTE9fmv8saNHcwr
svmAdwCBD9NgBlxJ18447CeDnKCx68Wr9WgFKwgc5397pv+y15yhwTQkDpP4CQZ/j0VJjz0BKGLv
uaDQreUhHXQayze0vwtvwSD6cZtEjbF/L8knpZE2n6N1XEiC6c1/mf7ruPO0oDTZzh1RZBO/xfUt
nuaz4U/1jGnLLQo7AGIiuNpb6PovJ5r9+fmPMHxmRHEBk1fXBMqbPDtYRKA+m7zrGUnp65qRSjye
GSp6Y8v3FF3pYojxMAcd7sI33isK67iixWcoaLqH6pu8rary4ol6BYB7YrJxQcQJb+Y3EeFwZGXJ
u98NPVKphThzuPcJPj28B6uZ//aM3jXpxy8NZ3ILXVnUhU66+oox6oZ7r5z8QS4vXtdjVmFwW0Ny
wWHABxaZHIi310XRzcksvmTMSjUcysiufo2hCaiJHt2YK/Ts9lyd+Sm+meMfgRdTSLhxF/FiImDQ
onwP92N5x2LdNNVUX/nM+hYvfLE19ckfK2vUYyRxo33Io1stRaPsNcWWlAUUEP2BQ9uDrzmCx+ZW
suy7tuXtOlqoLwHlKPaQyM7jYWhivymNTKcdA+dVxRUFqrjATc2RXVlAbFPVaIQ5PICcWM8iZl64
h20FLwTlwgNN1ek2EVxkXYC0yi+JWyJKBY1OE8xj1RGhAZ2VW+QQgLhuZRH+MpFJPd6QU+tAgpUe
kpqxOxffHfXAuvFiX9QGpqdXtHMtw39B1Tk/ZQi1tpkbQVEMXOjwBUxfQV76DeaLqTk9isATncBx
VepAStoYJiLaLWVTEH2aUWwB13Qandbe+WnVUUxK5VYXYQHv0vAFBxT8PjwtuiTmmqsmX+7K29Jj
bUVB58B6GpJ70VeoU36+gwTSoEXJn5pS25zJOBmE3A44bCKVAYgAwhz8n4lJwCP8meWfAdnfVoHg
sl6F7XxwSzlyz4M/wyUCle7S74oO06B3paFAwbcOxl46k/sGTNnIO/697FzktOMPYUgwagvgiaz/
T5V86Vo8JV6FjCkFoq2n3WAaS8nZr8F9xxoVe7Wf5AKEcFFjvJX7Ya28TsA3/G1l/35mqWVLYx2B
4gpDSGxPFZUNwJ4RlbOLnVhjtMcnMkc59jX8KNtyEsrT5/m2IpKT+OseDLJ1m4KYXyBTc95buBA5
kgkg1jc7T1PiF6ZY2SxOrk27US1/KfyxII35gyUTITLWcLHHR0+lnHx/a1hIlPchIFQkLYOJWDln
c+BTG99TLGgiFJy9+1v7aSSVHF/3IEaZLrosvu5qE0r1ekb1O9sy8vmicPiom1TVtWVoB3h7vIAy
LVm+F6Z32L7+r3WkSP/1MEaE7zFliET24F1x1Sge44YMj3YLZOMvI9/3T4MIyJcNC7wGwb06uIk+
1X6uiJNgf3IgR9Hst6rN+0n0cy9o5NjtKF2CqVAAUoInvrx1gldn5YRtzoMViyzLPImuCgIeD7LQ
vSW+A87AQOoq/HYB5QfivXhyiP6B0RxdaGrUmF9yXeuSTzIicPcxFf+wvsSIWEgI2gGorGIGeDN5
G6dT0sZzQwvIVKxlPFvqM8B8q+w+FP0iOAjyS6BtRGfQyURA4mnfk/E3vYuajAbb7iHUpGWNkR1o
MvfJE5XElT6MS6D286sIPrbSxns1VVitOmV/m+v19MkutY5mqP1SMaTAJDiy45yT/WgKb6HTTOox
nq2YxZQttHiYiWWI0uebOX/kTgJ2ICN2/7qf5b/XRcDw4+osDsspJVKUMRLy4B2w2L90/Yvr90vK
GKyr5muBHRnktokW1K3e8I18tXdfM2qjZh71bSy5qjbhhBO5EJmzi342jX8Ubr1x0BLn2TzzpbgM
qXr36CqpWZR3y6x0p2zcghXJBpbTHZ6QdVJEFw7a/JFIPwAQ8Y5RZgxZ8kM9KMnDWJkxAe9Bj2LF
MMXsl/yZt6UJW32WQNObQ2McV6jWs/M2VQ+Ut6a554+U1L4HHdH7HpzjadmQID0n5xslVAVMKrOd
pFv9ZJI5sYkgk8S4n8U4ffgQLLDvcOyA1aM9X1/o29UXd981TyMbq2XFP7R9M1kK4DwRJ3K0E3il
icAg7ISlp/jCq63rp8DwiRWUOINrX2WY3T+ViqXNbslqOeQAsU8rWLFrNH6JBmrznDXvIwmSr55y
BTXeGiCjlm+1xc9e6VRVppIizEQeozGTOPycdW9un9gPJybo3Cff0YdOYK5B0GLejd+VwcJNEC9d
fnT5IZ9Pp6ikbs8OSr6M6oFFWFMNHtTU+lEBZvQ8jKbI4XJsz9Cr+TgHWGHj1PM8PEz3LOdXsCox
HaLYn/UOb5dEstrS7MzyeY/D2eh7JKRKbum6cgZ8zLugSX2fzUt8oLJXI7sCwd+TkdICJRojnw91
tcGju7VIy577ZOzD5jrZSrySFQEgBB2LFjvDkKbtjT89lGru+vxKzdT8YirhXDL6vqX/pjokFaOS
ilUB5BX5smdtEB/sfayou/VtFhhFnA0AO5Qd5wjoPKlv1wTYIah8fetVEcf3G4h6n1rpioTWELVb
FEvtD6Aoq1eSPzURf+vpSmZHJp9K+wamIMsCzFbKRO2z0oFqfKMfAqJkX63ZVTCTDj+RdpD5i1vW
zHZoXJfvsxY+pFo9PulHXwUStrUNBSDrKBQ2r+F5ezC1rEVHW2yiE4U2WfUHfHMRoYtu9/a/soB2
+d64JAaYoDR3MqaCgwLafq45Ovkl+ldrNC5jgIIVuSJjE6R1fDdWx9t9PhBxQrIJabP2ska6Z7nm
+CYtIaRdzn63BBAKOteoLIOr6d0D5QBXSDsRkH0g6NfoFbIKaV627k7HKUL/2tNiviMC2DbVFmc6
F1HHTCqaDo4/9PPcW2kQ6GTqAOlpEFt/7If1d43wADc1hjlZRQ751XLA5VePpYCyrdT6+J9H1bfI
cyqQn7kvb7PPzgdWwFODB9CLivHqOc3lsM1f7T34rOZctOEKP0X4jYWARjhKFxXbuYIRc9Fi1wl/
bfY9emro292VVwM8yN2arufQsrG01Hx6rkIvct/faHjqP7WP4LLJskKWO6t0mYk9w4AbTR4TKKv/
L+84XmSBVog6qch93A/1AXMJu/7Rww5JOtrENfJLRIXpTJwgnpKph5VecOyKpFlRUTafjghgrvTw
PXd5gk8xKKF0DAHRp18iWEW5a4H0zylSzgsnHJgAbO+gOOW2goBRB6EWcmujzyQk4oaPLqNmS3Yd
pEfOyDBnVI11+dBehWbqLUt56trpvu6AGjPLutixvTErJ9kzj1mnc//LfBF9/HhlHAR/FwEWc1ah
skcwWBxjvYz/6faAv5TArcvdBUPMJGI28KpPV+WmlndWOzUG8bQgnNXICYaqd/FxvSGJXVlo1Ega
dmaRxXt0DKcBcGvg9FdjKI0nneBBFcs1AFTG6csKXbYdwrPzakFk0x0M6EYSfJJXTfXmwIu9dqA0
8IDv1uecXMx37gbjVk7/yPiL6HInOpDwRiEdOJG7nmPuN1rutkaLx/BZ6N0kqjk94TIAVol2yvni
VTw96f0XzTXsjmzM5eq814zxO0myvW1BFlOMAwq7My/nh22e6Zzbc7UYvxz7CkJZIM4fEwGgfNnP
IH1T17FGrpzsoDwghiXDXFFPEIJDHB5mjPw26RUPx3XdpG+Kq3q7PW8Vvppz16KwT9SfUE2cvytD
wBEAYgm1shBOBUhoGK5MHgEpuAlqgdwmdzX65AaRdv6sMjAdrAtBzB/H0UsFS63I7PCBv+ZZfLnc
6BGnH7Rq6O+Lqc7I0t1hg+GSIkGfSqKSjipCkXTU3iDChRAwynyLn4q+x7quyNe21LZy3/yEjWLJ
u/oVo8A4jefmmV69TO3g0Z1EZb1uSVJ4gr6CH5Deej6h8bCuz1W2v9k+XL+qttu9SsYoRAatEIvv
8JCdSab2nuHPOZu00VxmhH/OzqvCKriD93L3KFBzyYka9f3yS+HPC64gJBN/NhWIAAFkpSqVY7/r
DhuzdGeRmGizHLub8iALipj7vRN1ky/IH/nswOwXgq0fA/1Kih9jOmRYvDntzKU83YPZs76zLNUT
a7yAsHZiw0dJh8kC2c7dCePeRkw0y1F/scFpVqRpsFYZ/L2eU5EtiF/4RjjiI0gFzavM40kV1S2e
XEoW8CztY7GrBw5xRhqy83BUmmKiCrZyOQ+MKQDN8AFgQHTe2NirEel9/dPhHUFN+6gnxvFNESeu
TS7QZjqlQUwkGKA4/pdnFrrv3FQpfLImqJdwNASpXO30OGSoiSNncexip1x17d2UkWw6pTnAB1zQ
28d4btxva841JULhEKnrwGHoSbov/p5nwwEPAHzk9IjFie5oeovYX+bzdqV2JUhemEsB4W/R0xo5
Gd5NOo2pdflJcx9uiFqaBOWqKMHPPXHTB4MVgwwIwTRy00/k+9CwKXMIZdMzsuNton0Dl01vAHJG
3vkyR50rVJicDkFoRU3TU0Y0vHPYBlxi0MJZ0c1FqZZLlSh4n3WZoAcVy8WTz07m41xroc2D3z0W
0VRD3xDMvgzXicbXCjkCvURb2cxYFAp8Uv1KFnCeC01QZjF7xJP3DLzYJu0csj5h40UeS3RwJ0d8
M9AtQdFy6xALAyEyikwPsBbiuv/ImN6rgOgohr9Iv6IXY2bseQJoyRNuFdpYH9U47XlUsrjApyda
gRJ1DHENowAEUk0q4stIOtjUcPBqhWQR8tJk/yinFWAy1DKVJdQ+Dzu3i7WpvwFBYfARManYKPd7
t2L8gNqB8TX1lfGG/Bn0PHmg4mTeI6U+ZdEGgztgWgnvLb1yTlX1VfLCC9IC6FiHnelGndseENBR
d9vxQpVXiggBeF+mQVeAZESRaiIehKLvM+5ERS+hNHl8j7Fa4M01ojtpRuOLxQO+U49mK7O81iiQ
0dMg5tHNZT1RcAmCqinma5lmazLEkSsWYE0B/0VYK1dsri70A3p2pKtplJLVfAbmI/sR8umU8LPT
WRLenQlAtuCWdaMUoabmtACL4VpiCPuZTQFQ5w7rQfFYB9xLMQ+Ov/1254M878twZH2Dy3RZ5ShU
iKi8hsqiz6wYAIboCbzac92REBl0pNDZIb+uhL9+haCjE9kOEP1YxrPccI4qvgp+YNa+bEHwI5zC
JJEyxXht9i7fPRKXlZEfKxzVDvtpXa7AvOtJJxpWAcMSjKYQisvidlthpr50BEgZzun0bjW1uWtV
NtjTqpuNj4hFvYwu9oPRkgzZKq73qB3x0hJELzFA1XPyjbqmx30AQGUrYTLzxJBs9Cl8MBWjndL/
DtCqL0FmuR6Mtl2CmKTgBnDwSuZVU0VQ5/odoq+/dtISv6KWMR3iXtBFgjA/AHZ/WNl4B1aqtjDb
9vTdcPA1p1drRkeE94Vdt+DUuqQhwa4B72jF7UZiUnF0xNWz0OmtTJyJ+8jbXbQ2bZDy1AfiMZId
jrN+QH07yFc6dEvLUp6VKQwtC4sdtlyqz48SAMoZwHJcv7eTBZ+R4d38DE7RWGHfaLZf7Fpwl17D
EaJX7zuMV8sFkc9CRh3z36ZlhmJjYMy5axCgxXkXoxi3mJUw7JRxxjgxVW9GYL2DmdjazISmMV6Y
zXJQ+xpnP8RnrxO23hmRQrZmlj3VME/KkXMIsajWAL++g8fe/2/L9vjqNyP/H+v+y2BIKk+Zf2W2
uBCLBVYlm2x3OtoH3VVk4JvcZstDWsqBfnc03JlonKMlrmdAGJiRYWhANOACYVbx+mAoRm2zWCoh
7dugLjV+/qzhRtpdws3rWpOqPPC5j2Ls7JelMPOyLqgN7r8b4c/OpdU08n8+ypZ4NpZIKIjN+BQs
DN2GvGeFj2HNrq3eULKhyCveXIKAKik7wWxkGnBw15Yw+jF58I7EiNjRarabSJHNNosoIJ2faWkp
MBmYsW/Gz4ooQsnjFhAWDp3F6gMoZqBKvAs/3N9C9pjP6k87Z2h1B9wc3olI/B9gHV17/vR+tc2D
0Xqt9+a7em1Gf8/c1lpmc6DCFHjeP7b3l6l16gMup9sAML5ynJuqBNQ7AKY0C7AS47EoxnZoQfy8
30diBQQU7oIev+411Op968ll0gbUcRHsjIMEB725iVGm6flVh0CpG9DzePieRfCE1qFZ425k/tsv
Hi7ohlmdyPSRJE6/KMu8GvMtClik9m432OMwuQRoiibMv5IKYaQxsIHtfFOBAHyC2RO+BG2Df2TW
ys6ij4NuijwbF35AS1m7HFRECuKrqneypJu/j4QZEcuTabLLsCrbjzKRL0UibsdCMV9DIOZatOgb
0UVFEX/h7KEILPkatikGjM3iB7ZrY+HtPF40WOcdRfh6I6RsVqyCZ6nB47ErHb0ZtPzg3KUCe3Jd
3wCl09sAquLfJulyF+WOa56i01WhQ+vGVF5lDq36eWceYsUMHq72t38lIdC+tPhhncrDWc4MCaoq
mrsfoI46lTsiJhITb9n92W8D4TCwgvrQ+eUVp4nLPHOy3B4JkG7u5AIHbo2ertQp+r9tjXOpi4nE
UCvjBHx4+h6N1sMQwcfkIH4hB9jk29U0Gt+yZDvTNMvYnAGkLpP46hm/y0bAepmzRwaibsTySDgz
1TQsXS+c4F8lQ0/6LT/WnprUaxVZshU74G4vUqb5atQy4hhWxXWg6DFuvnfW0EwDSZGwqKHLTvqN
01J/0v4KeA4D+P2Ch5ziH1chrudTgf8ByWh9aqX9Nwy3SliYpy86zWY1UzkEjoYlzBMwLyBeEJtA
R3SndyDB4G8Iq1LONjkuDRQFYXYYP4UTXh22zgDmXHTyjONFpT0mEDcwNxVWL98whCNoqIheLYbk
G9PVP8n0y/fc6I8TwBs8SNiGUhOQPo6fSl+RIzvqLxMUuff7sope+JSLf+3y0Wfq0N4gZ9aYykKO
Ez+h0+zaxaV2EbzXYuZl6JrNUSn5xGmDXIYZBo0tyQ3zt9A0tg1x6is6vYlZSL9896xUn8psQFCL
lw773Yd8yFAVKiwrLCYEd3zXB7TyNIeUq5x2CvMKdPKo+wxBLlgti/zwERle1zqc8G3Xdj/FSgsp
xxP5iZMGLffICP1me/PsUYq9i0mbCih5QAYoFtRQtEWIE9YulItlrkSOGnsVH2Yj+xXgxihLh91w
QDUwfOCmSebB2NhfH1tlPfBtjsjEdjXPxh4e4BvHZi9kSbWg4nbupqu++yoH/uW3j8FWNITP8RSW
BSNmFoaBx33avTqQT/rd26pBqMuKghQla/C1ejhtXcc+kpskweGhjk3fU+5njx3qhiCbdBuATte1
eJSFvCVe5bix2s8ZdbuyzF8hZVKnsTZSKU/Sfp4NQWCxwhPYUu44genlXzP2vcOvSPJMzVAo9kgF
1LvWgxVsEdboKSaGbxnrYIbnx/Wm+1t7/H8tTqbWiUsiHQ0blrzBPnOApZPhHdujNnu7psTVp0O8
L1Ne6FxPuORDCDctxNGhc7XESTc8hFZTwnzCsAcz4BnlM8rBuNvHYZ60taRZ/yblFRo7wVc2IaWk
2jzDqLXxEglsoU6mBNbUl8rB/wLBQkvU7KnS9K4/EuZSZTDPWr0gPMLkiJa6bVvyrTF4yXD7/zu/
cIOh0GmKybBYMJQt/dfoFRa4IeOzY8i3w2ooEvy3cSJCeRjwPKrKrXRoMT2GhOHNZsOWSLEScJGk
lMR2W5H70NHN03xCNoOPbe8H7IM/xhjM0wQjUwmtCqgXwuUStXCkMwFTGUpfUq0gkDrQZfvPfGxx
hmCp4YnzCKpSq7zvmB8i0frzpZCY0+6LvWeZdWw02RzM878onI9tUgDiog2vEcw5gY5jPImf6/oV
M5vCCP2lkrp5t8CauXd3nHTPynRmlJg0oNFIGbyD3VOrxch0a5ux5HMwDf344vdlOWeIJtofrQa+
sh2fNAultMYWj5tgKX8oI+nPsawX9RXqL+W8rq59NxiMeuW2ObkBFV4ms1x3JYUe4VeRTm0XsXRt
dhFM6gAt6mTLzOEpuYMUYHLKe0WBcBYKJ3rre9AopAeatjfJUu40TB+rxgCgT9loiUk9AFsugHku
m+hPdkma4wdQbi1UAlD1qHMoqa+kJX9LDQJzMJ3fvl2BJKndDH/vHWhn5HoSmYajp2txbQmwe9Lt
RRO58YtizKKleoTUIYYm3oeQ/FTYhLFI9/XP9vsgJEDC3yK+XASKrcW3OWgCh9E30Z5uBmSAm6ls
HqEMYwwwjlLoqneQrPqyK55sudNYE7w7sGM/8pLcNqgpKQw+vkGMl0B0ce5Ago3LzZX4KoaVr0EA
d3GuO143WvaxupTpg95aqyt/1APGKXxTFREF7ygRM0Y2l31A7+gu7jI6Hz24O6bVGPbsZe3wbbtO
Y413WFNGZs+Y6iiXEfxiQwXhLGBIoSRAUDdTv+E/j169ZGvlDMq+1/VMEg8Vve5qoe15lttxxbB+
uUsB8KwNR0Y5eYR1F5gaQdIeiYicOsobgtzwwOqZLItBGElHL4OBBfxmqYXYr6/hlFfery5NQPMi
zD9iZKREJD1cbkYx2CG41SV+9V6Qj88/vUSPJMFxPAcvAVSyZ1oxhlTE0lYajHVHsBvNBM4joLHW
svbIX19pGy39vVByBlgA4nRJCqyHzIABrJBq32RV3Z/jExIpamBSdZz0XT8j6GS7CvHvuSo2oMbi
XD4ZZN0kdDyj2OxbMqX4XyDw+TRsub+JnSF4o6ssXRs5qmvpu2pVzjorOFjj/w2sdEULs+m7yo8n
CWDcjbN/1+j6QvCgefs2bxV7q87NMplKAkoZBqRjPSB/dgfxJi7hGF8MGPc2bZsr1IrSwhlx8pvo
WsPXmS3XZU4IlFwPvcQMWpsmbobj28Bx5cVW9Ee/09/+rDGceG1b6JaZ0kHiugCnkVxsRkZUluZc
v2BpawBPHqtce4DFMSV29GYrk+5ccZrRwXhAb7WdJokBs6Vj26HM2/xS6ADBd234C/+7eUQxpVyz
9Xy9T649Wr+wh9eixswKWjR0ZCYQmj/b05Y9dQyC7YpDuZ2Q1LpFUBEySY8aALA/jC+HTzOK3lN/
pZygonBu4vu6xQaiN/GqGX0TaqVrxxnjpdky/IKr7R3haAvKESqz2hvfYYgjp24hng1KGQEDJ1Dh
4PTZBj4rf1E23qBCdXQxttIDnHctP5TMi8uWSFbSEvXjzx07YAJG7upizkai4qPy83sjxM+tt7tw
sairPS4C4SNPZfMiAxUNaPu20O+EQ1ReFygg752w1yEIpEJehG7kZcSzhsONARy8paG3auEPw/gP
oeFjyyEsAGoKxi/LyVIqKA6uUZ8ax7d9mEsCmwvCv3MHYyZtcmacfGmNifLJIrnNUCZkE29CFrT+
GAFFrcUtiqqT45W0+Ga1YFHWpfCNMwNCPeQ/wbA1eH4eCkm2wbiC2sa3yrtXa+7X6uzRVzJYb94V
pBkf6N6KxYSnvAdhU2vaarCCRZVJ15cx9+vDGQ0JkTcdfKWpDR67wl9WfWukjYkZccNsCojwrXYF
nYVr/Onlxjl5t1N3yAc6AebOTGyGcZJmscwqukoM0bZ3kymnS1U4aNsizJnEYhJCV2CEj6aiIxW2
wOdNYBF4HNeQW6yjyLZ4+/M2MdtyzeqzUvj8wOdrHLS0pIhosfgRRlDOhOrj4lTNNCap+nQz1nIM
ZgG4yu1RoV2HuSZSIcMH86HmqtX4n6/+OXzgZqqubtxxJHYqcTdkzB9pILuaK+MFNEmRsKVxcmTP
N3SQ7FbvDvURoE6PZN9Bw7QMDjCijyO/XYzVtibnmPS7SvSDOY6/tkgNKGrJF0FhQNf4P0kesYrz
G+7J6EX5HVR3ifsr3zCabcmt3rdrZACH8D/s2M5ehJfPV9bAlEjbIx3D6JS6WJkolfYvPsfsk1ih
ZG8pJW6MD0V4GAnJ65PKfpwefpKgVfqEvWp86gvxtCjeFzuIGD5pNyyiSVhs36n2mVltBlLZ10MM
mqvzdRdXT5utqY6MA43bx/6jMKETmbD1BTEXsniAWGKEE7e9wdOyVbG/DJFyfIPgJG9PwYQB6SiF
dOUdpQQl7n9DjaHJufbLmjg5+daEFcv+Y4wEJE7DaLLZatUl8wDb9sYf6MrZcYg9GHBtu+9SgmAg
pZzdBNZcxW5shh5x+72J7zSJ4W7+ML9hUlwOVt7AIDxmsH8HMUaBcqDwctwHMkIXHPTV8Walkq2S
d6xuBRnSeiOC4NBpFMabU7qc1Q8c5gtcwTkFYWuX3MbirlkJNaJRWfyr9V/t2vtGMLpG7/pNgO14
Gm7CnPGoZu8WI/MdFtWNw9iYJPRBfklUY/Ehhq4X4Lks28JRNTYchF65hwT0TaFaBuCAMnfbFEnk
XjAqPlT8WtmUtE5CkagK5FhpbE5jDLxT3Efsv+n7L909etp5CkBwtM2rmcp+WFfshT8Wep1qrTKd
Y9AL4BL3oJT39AssjyLxzzxw3mMpUklsKJiid74rlFEkYvUzwcTCKXAG/X5I2XdUVa+hawPCWn33
Qm3czdjqICjS4oXngX3VWhRHTSVsrD9SgbvtcxzFtoTR5CXrehjbE6dRhYkzad59pU5jC0/sTUzx
wkKs6/8914knO9I/oSy2Jo48TF0Ooqs30ZYShHXJR+3bptTYk7McUGvWNaFzHtj7a/Ol6T8ipy98
n9f/vJMvPa9AdV2HIbMAfM8nvQHfrtYDBgWielAchFu6qcReXJKgLGaFbOzPZqKcH5E8DJGmHXVu
20Ea/mYYUdOEifmksUsJ+G8FnaJYsHMlXKjm1IK/SKPnLGNsy1C3g/0BrLmhhPeFomxp6suvcexo
PgZ8nxVHfWYB1hDp7eg/wKtIb8FfjDvAVcldQMfNIypAVcfn2ZQ7eDoaMaZ0mh+vIoe3MdWnYiOY
Cf/D0yN/UMzrwdZVpm1ujbia+3u5xT1W+LaIBY4IuO/44WuxBw8WAStSGaN5ux1CVPLoqv8KXWot
z0BsDLGpGKrM4cks+YBnRz4pY30q1z2aSThv4NJta1pq7JJoyDJJYMYbqfc8jf3ONwoc5WktQ2Bl
M+G0VXiRybcDu8UsSnTfwwsE4iLuoUBxDt35BT3vvU9c8vpMFb17IUUchs3rdWu0gXhIKweyVdlZ
fl3+5ZW3wRdC3ugEiIZ36N6MnwBJs9NYMYhpENrD/+ghb9QF/moQlh1XTGATtXOsAvKQcogNC9p5
g6SKea1iXG7Xm1E8KYr8Q44gWuGskcT3yT0GdrqmHFx8HQj7qWf9weoR4FBmqAAaiNrZdbZGDuSu
2FcxeF4d61TzA3BbVQGweDluMc5LDs3ZenEGD9/hFkZU7Q4sKZk73qxhcARQcdcYxGp18MJZqB2J
tGBwHjViMbp8SxmTTHgTLHIEl6bbcWuW3YKCluGEyzLBNe8kpaNkjdQPSOyEY4oeHM/MjdAInZtk
tAdWRg9VGwlDt88D/S4RqxAyu6vqNxEB5J9ir2+eL8u9rO9Umm0Jz8SEetY+PMwcp3HUXRNXkHuG
MMasDnQv+FeIjyZXqOulXzCc80LAupvh94nfUA5VaTBaP1IT3UREYcXj2yzZQaoo445oprUnrcB/
te2TpLRmjicZU2e6WBbPEQtXF4qZRUkYwQ+oV1O7TYd6Q3744JQj36QoPNNvO9aNp89hICjGnBDs
rTNR7cYcxwMPJ0jrdg/N4xw/ZohU+R8gaXPOQgq+RHykT/lklxf2oQzPHYCCv5bdp3EnVJXtbyor
4iYxbN7h6X+adO/tP2vItp5AJDmgTAp8ytMiIIibN5qTK47Wnp1fJiOLuDZ2Lg+nBMdOHVx2kJX6
JyCiAcDAmP+TnpWqxBZOpsdKtsTTvCRZI1dOJYAEjwum/awEEG+r0Ti4kaaFy8DhKQyUxsxh4Mgg
U283eUsU4z3miOR3u2BFqC33t/nsT4TyHIKdoAk4hpARp4dZDDROBk4EvKhyPS9LQIK99bZqZgmw
sr1KPddeU3TKKaSSkvdd8Jkwj6ru042d/5L9ZagMXUVIeJ5uXblA4ITyMW0nLwkaSE9BU/ni4yXU
ig//ImhuP7mxm7+D1NYGbF4qRyKSTblTzzCuU9BAC65mRLx6bKAIK7MJMLeOqmb9ZiNWVtOUri2c
ZgS8Qk9hKHCiaXCIhYG2oN5pCyJGkDnVB59YXsBCqLKmyIC5/RlLkg/cbCQ/3QyPWntnL4erYDA6
6IJx2UKqfnmR1W9SiH/JGlUr3asb3VN0j7B9fyL2XGU0dwIGnMvEjdrHIQK2PyVq7N4XjBlvn8p3
LdDbpbSvGHhovX/LkuhDBITdsEO03/UKiHoiDzGDiAGnveX2GjzRbDWrkZOWDoxbaaIfKyV8CLtq
tKkxz79dqPMxyoOcwzzJwh7jOWUmVnYUAhoybhpKAiPZ6YhLG0Q5Pd8BLz8mfweXORd9PMexs+/A
eipC9cWODkq+SqBdtUMmN/DNovMiBc5BE3CnHBy35ZcCW4IDhsizime2L8iyxssMEqLb+krz56mO
7OU/wBjme8EqieFk5BuEHbczTOzaVGBQxGUwh+tLl5v7m2P3cmkC41BgECf8sZe0Kgb+zgCpv9bv
dFA5YiMtpj+Lh6Vp3wgWKN7a2wl660vGWpQVU2N/vOCmfr6U5T3lYv3ZXDEak5xN4nD+BtWE8pol
GXfIdHjXMtc9204oxz1307NN4UkIwkmx7dFnnVDQKIhY75wWW+vKyvUp8w4Tt1sF7We+7HnaMWaX
Evi3WjyRQ0AVs4WZMN61Wfr8e/Q0Eqb0CluJ3cTrRJkV+4F5P9qKbqH4X959XCCgOk1Itf0NaH+0
SCwfu/u2wShL3ZeAYGKYcBQZicXD4KIDXB8ru8DE1uVwfdHCc4Al88FOhKe7RP+GiHw6nvrFh7MF
pyYBcCv9TkstCslpAnlFIedMjVxfQWmegzWbSBH0uVB7d++RnCgujYfIm2sANzp5ZAJXfiZWSV2w
vUiUER87ZuaLQhxtnWa+JjsD8U9RwuuLoDKXbZeEWu311sS6fkDmmQ8Qy4ZhSpYz6WePvNZTdBtb
JoSi23PFUT49MF/50AS9ILNlx+hemantuV1Zbd3/vUqdFMoQl3IV37k6elzhbMyHt22DJRoI9Dmq
FrTzS22IEM4lSnBly1Q4hXxtON/GHge17HmbFU5mE9GGqsRw8B3xh5Coavx+WECm5s17410HpSJI
8hOfRnzHoThqZSH+0E6dosabcZuJm/cg9QU3PXT7QxD0PJIrCKt7kfP3f9OoEHMvGT1aX8GhZV7C
LrfoKH4cdhjW4/qQ3/nLrtkLQfiBgKJQYCaIL+6Z1hNqurRG8s2LWoY4l/O1z4+vLfK6FLSZKRFT
K/ArdnUYk+qy/HfFGoj9Q78CWWF8dnUm8zTvcLofUOmsncw2xdiRv91GNZuZv4lYolYygupOtRGV
fhQZUh19j/oirJu0EuWxa/JVHVqmqZ5g3TiC9MmMdz5cmemsU99VFTWFnWXK80LQvGakalEpatwl
iS9bDlrKj3u51UNQEvNWf54wrgSuvp1sqYS1Buf9Ufx1pw7ZsHdsYF9gDPK0yhUV1nVCSiP9mXk3
tuX1Zg14K9++QTw86sNRk4s33lcyAENtwiOlJ8MucsRi3SHqtQOwSEDAtCeXxSjy4E23zxrvPVAf
HfauKdk3HvdbSnHb+JL8egAOy5Fi8r+lqFg7x55hHdc+jzeSpeT7937ZpnYyL1Txr+lZNTS3k6Za
Ii+YSug+j2bnQKce89aO0MG+P41XpzJ2YACCd4c7cexzBvMfOar4hxH7QN2UHjRF391YdEu+kbEx
shRZqt8Q9Hp7AORsevu8dpBPkZmGMXYNZzZD1c/kfHGsDLTmwMPEpQoEedi9Vm6qDIa6ypOxYrqH
dFbjKdGQMHg7hG5/nbZuCtnDueZ7DEkWzBcAmeyN5z8kLSR6gkltEeEi5VaaBWHq3ba6WcVO5Hdm
xJTzma/X32m7BuE2+4h2hJNhDke1+nf49I4wVRP5Z7CvCytgpDAAUULSGN11LSR+yB2sjs0XjBXM
+Xm+HoOD++gNXYHnWtOOuWb3uj461i19//65T+Nky93nH4057e8WYl3miszEN4/EuRJf3JsfiL0m
WJS4cGJ2l++Rh5DzSaS6wmS+J1bbUx3NLdlPPmkJBob92DIVq5+mCP5Vbz1EPzGD/jnAAlm0vXbZ
ORPFzXwQ4n3SZQ0lZi/Xa0YLIYDdhLA4HjSrvMRAYhfjZA3jgV2AHN6/6a/o4aDYDXE0QE96hUU2
wdezFWUnu1146E/NNensFkCAgfu2o8hiuICEnaOssZLiKHttngaMsFvIfA8GAMZCiEANxH8DgEf0
3+773i5QG4xGU9QzsS4fFBaDsvJf9YRrDuOEUSstrS4gAIu4mi4sHEyRq8JUTjWvlBZcVbfUD66/
dGObFsbsqvhqYGp8cjoUldCSAk3BZtWCi+pKhXyoH8AVorGtzi0+YOQ5KkpLjJ48T6HWrKz8KyyU
gn4qnb90yDOsEWCPVadgNT4gDnNKFs/7Kx61K5X5NixA6TQwDeQKEWXkOqXdSKnY4iOFJQRaiIvW
SdpS2907D62c9EjRV7JNml8ovM6ugkHumy160EKpjGpFpkeAj1BzGpRocErs9WYH42BgcPofQaCf
4oIEKQ+QMhaHDZZlqYaSr5+Oypm3Kl1745z88Z6ZEPk0aIwj3J++k/pmNjNHMIHWxP8HRGXOj7a9
X+aCxuwWhQ1tI+dCJpgZK0/qJEbHovm884qRg39FUoP8FdjCYFxm2P3JdNHhjhF0b6RRMboPwYvd
QsHflKrtLrsvPUH+LgZ4dKW+be8xcJ+ZvAgB6W9YaEOvlqgcfl15X3KW9/PJa7X2mIlI++mStJBf
5H3JwwmvWqEJt8LflgfSkhqnJuDREopggZKBCcN4tVYq5DlZB7Vqe+r1Ka11y9w6p+QL5F5QL0tf
Wj3ZZBcGKuznHBIj+4czACivB/tTFNyLpTBPB9UUBiRZJOxZLpk3VMF1FrDNSVI9Fo2VWppy7YHD
9AC/A5CSX5Xe3yI9WjnCcA+7mXsDgLO2uQ1B5wgNLyv+MSbPN1VQdxPWLxcILag+zTXOXwpNZNKz
o8MsOmbYaG/PAHaV5L973QR9hiWNg2J0GqEXst10HwvySlwp+r/S2ag8lLZE1+parQHDalOLC/TV
EKQwPrzONvpyxQylk+l9sZX6IBMM5xeRE8sijw0fUEN+X3E4k1T3GFGssiTjotWSRAcQjeWS+eyH
zhJ+CVzsb1vWzDtM8ABSQjilNla2X9a2HmR8v/vuuzMK8ZaFYAAYyNjTSAc+etd7Tb8bzF5STljK
XXMMRW7un2d6wNL66gpzdU8M1lE7ao0kWuAPWk8LBeTznrKFdSEqCylz4xvtBvtol7ZfcT3+yO4l
2Impbrmdz3h610+1OgdDwaqDwMejnNmc8UWphxeD1WlC6IZTQuHfkktQeJoi7JM5CxZpo67daGnN
fecR2gERDdYligS05Rvt4wi3iQuZs772uAiUuHocOutSTosZslcbBYNel7Cji1bK5/UtOz+PUXKK
5DEmKzNkbVFiIbdBjmVIiCO7f7c0AavBdZamKJ5mV+cd9od38GHfLBa9yh5jjlnLjyU1HT0AgUbG
Yrvh3Nu7/fpk1ET5qael9PR7AWfgS0RolHIUOqQ2e4hunlR8Hq8R057JlxExEs5/PQvKglhFIlHD
6R4cVDJ/Tb5HXAyMgvxgVqLRb+Jjayc4Ao70F/nIys+BmC2zp3+alNpymOD/H7ox/IMUF2OhTVWd
3AfgyKJuEM3JpNoldtjbPjVJ0TAeykibw1q1diCLIOAgK8mF01A0hRx9vzMUnzd1aIBuN7poYJSX
roCdj6dsN3v6+bBr5MGD/pBLOtkjGGXxE5iGf4BjFDVKLl0rheqLcPKXyg1lJ+0/K4pBQqafOIAL
nVGxjp2V3f355Qfm7mJOTJNQ9Mk3ieCtVSsD1nLMfxhNFMupUrMy/OR6Hq+cz8Y3RVltAY3iJO+K
z8ntsSBChzirjaVa962eUYkyVXapCC0LwNWHyBbAw/N4TfsdZb6D+36M3y7fVinjIlbfZjX5rFaF
hbWYfH894GJ0mxpAa+Q7EkXNHVkNJpzi1wh0gpfbACPTNKZhWmpR5HfXT356LEQpOusmGg8RRc2Z
7iLB54kza9XkUBMMyRKXRua1Rj1rPVgx3J8wSq4Y2HIni2zDhJJ4St1OrZQNsRkywqC8Po1t3XEB
IzsUcl7xMogCv1fTzI8f1RqRfAdzRfol+TZ96MDjAgaopm4dZjKjmrq8AcMpcNXliXLzZb82LP/W
jCS6KcxauncaWYwPQO/j2FzBIILWuZ0vhUqONAcYmmb2dWjSy0IpLitU1ss1JDSGk3vPR4ZpDoGY
emEuSahylkIXr7z6j0HmCphHEESlVebi4RkKlDVxVbDL85wJvvfmkxZeDZaZVwQOVX4yoi0p8O/O
ABjl6MZrhmSj3ivkmzCBhWaSjsYtr89WmMtk3FmgOxLJtM3Fj4AV6tWGsm9A4JfBkIofRQfhvO6r
aKjRsVI0X0efQ7Yj7GgPYjEs665njBbgisL+pNp3n+e3KjVF94n8x0gH/X0jn+kLcyvW8PJX4BLL
yX9B0rHxxlVbvn3iV8NuaHZU47uq+1+H07lq0ukB3nlB0E4AWq6F7wn5NAFqJ0f5z6f5a3ujwCK+
fTSsd3vpRz1+LVE6J3Ak/YL09XQkaV33QdyitVLQ63JuE8+c0yLOVbbRk/wJx8/n4AUje2Z7A2g7
G2cSXfUhJnwcO5NsYyWeiCn+IXzGwCBFH+MdhAB0aXM4elyPpeQ0DWoFL3KvmAarPz/iiPUrclk8
aUCkQSMjCKE+dutnvxGUxx2Vd8jzarVeq0+1jFjxWDIaLFYrDlb01HyN+FCrlv6ZEeDjqy+FB939
jp9LsfRUy8KO7Qoleczdj+BNR3NtevD1w5Ze+KrBlr4dCyDN2G61eaIOuphzaY2O5hxtHTT2U8by
Ehw8pPLlHAs92osBk1uClUgoSy5T0uCOGLgu6PTzPiwdI+dHiSVW0pjdmZmeTUGZt0MQS7bLBbRw
MOIiNfNxDwC6m6HN6wDSgu4gQw50oU3ecWlrLS9kKUWh00IzEtVA3o73vRaFij+XfiT+SKg0IpTH
BFP+1xSZcWRjTzhekPmR+lOI8YpYF5Jp0Asc+s5scl8QR7m3nzAG1x98uQqdBWPSuR7Z+xGE3E6s
WJ4lgPSbIqax6NmyWt9Z+xNwUFs5P3mPNDJW5WhG4o8epl/C17N8qEp/k/k02iUvJLLBOcaqG2r+
tmCKZ0ICvrLiKL2zv7RwK2LFnRSHUta+GiUTjrNzSldOlyFOHtPCCnNhcrfbt5MR1QExKLLPNQhs
D2o4M3R43EsGcBuzakOlU17nJB+hp1Uha1YWBFlDDbJlpR/yaZH+jC/oNlgWqi6BWizDByoFapmN
Qx4JCzJ1DGge0mjA+VvB4A59RPxwyuxIC6QSjbtX/GixwXH2aMHsukX3ParbBCbtAACVz859FCBO
QFq2BKFjSdVpJNdGjYtcRzjixwVesIQ0ZbFN4QooyH3uTKzgtU31OWCG0wLsWnm9l59lMjSToU6H
fKK869Q6XSzuhxEXD99uPq6a93zmkjEE7I2kuRK0592dXrSNdmm+EU+z+Rp8Idsj4zNdgRIzYbRL
KdSWWelVvlEpeZq7s91TEJRLXma8B8cij657oRNNzHQHHSzf3gZU000oJ0gvQs11vRdtEFcL3NzQ
0Gph1073b13he6WiLllH71VpwPDyK18FjJYbXEEJJm1Y6FrufhPcvdPgGT+Pod4QnY9Ei3/E617c
Gc6aXmrvL4pSdSghFS7JjzUEaQg9xLc/syihY5uOiOkDwpQ7Q1RMqdgwoN3f765fvjBzwI5ZDRtF
LMskoxqvXhUIi1TrJxcl6iODzoSD9DIJVmMN/jU4e37qgR9gMevB4voQdg9MPMWEaPA+2Ed1ldpq
yQ1McHj511JUiE/2OfHfCPXiQBq0qdqsg+Np//AdVBLIkTF3meily8Xm4XJoxvv3S05qqFmhMM0u
+MFyfb2tfNuPUHFuN+m35lAIQ+1ic/mR1HbwNIW9ckzOQzf2SqhRxL+BJsSBRnFpFKjzHi1QXpVo
IMaOOOHtr6Y83oxhxGJ/JV6Z3DQ7Qkvp5SS85HfC7lbXDrjjzpki9BJbECsMIiz19Do3eYuwMGSB
Ut+g4Ny1OtQZ+DiRNcLjg6+pTVum+xNNTNgAGZlx19BipRDwf8fCGYB4BL+XJZSZhLSOIO6dFMQG
n2ZcYe9q1meCax8iUQA49El2e/6ylF+lck7BwnntsHGm+CPCeSxYh0fdop8yXgjJ12XyzK+HkZSg
teoSd3rNaIVxtVZ1cm3Y+kO3JXhs8NDN6lFqr+dgcpn7QUTe5bVLGu9Ghc4WfvX7PSO1nAHflQHU
rPGxRi/NVHehVbKadq4QheI6vX0atiz8W3f1ccR3RvPbsaEJbSFIodBApfQj9ivIcbORZBirNxu8
2K+tTaS/pdxVvv76dlT5o3P0xsiffex12Cn0l7fyZgmFAcvx4eH34SQn/8ZHkr1OfOYHdBxSiigS
yaXXP9CXvuqZHokB7zRHxVaO0v2ks2KPLYU5AJ47Tyvy3XkwYmrw54ayfY8MFayrAw7l/2uxQ6VS
/B0562sH3lvRqO+CcYqSmY67lQTXrEX/4a0JQpK5ZcvaMH+W/PUeYSHvPCHeGzo86pzVJcXZLfkm
nVPUSNIfIgzvKTJhRr8lxnMGPOB9vHuA2vMOlNp6cCJn0JXerzcvgJiVra+FAP9dXcK6ZLvUFt04
nvD+3E8k1GhhHYdmuSTdTRBpLdTcbTA886tbn2DxG6sDSWFNzpC3nqUb/8QfUB81FWDwS4ZLv9/f
Dx3wt4oAMU5qyC0HGpaW6zYbEqqxqSayXknBwiWHI3W8ffW7QaTrVcg8FmQjUJg2Uwwz/j3rDvky
UrrxRqFFTfAVNSUwuzF5lfugzXTuYpgQqSYoQjZsh9dyw3N3mPDIiDFTbI3PwPQ7RTYX2w3z3/BM
NXkyJPuCFvXJgbXBlpKsRCb7kczqU+pHvbQpvrOWRMt+VgPwRjOX9wiU7awwnPYsP9URpllS/338
O2OIZMUvE6JvV0PSw4CJMeYpa/ZeUndmawMproaPBXX+Q9WvXWZylDTHBQEgnhP8a8vvB4Tnrhx7
pHuPmImW9CVFNLi5TbAGi8RgjvQnTwHH7pdIwNg5XGozHuFQKrlyQs8IS0H6MONBHZT2t3TLS477
tfpRMVCPxHE6ihMXAnLs8OcNLe6flB8c0pe/60zukP5UGXswNl8Fulz+5rmEutVS6+KHriGXVCsH
4Oh0bKiKGpRxPYzXR2+c6DZ3jcTkWQEzvXqXPQ0C1bNvXBc6XBTGe7M5R7mZc0N8IpKv9JTi7H+0
OymCGYZm0fstEehUUr2sB4yOaCovGfq3zBx/hyxz0DEHV8AzmrOXFGUw8aDfHxx73O3n8hSpCYUj
MqPUTLfH3NrDRlRx9NoNby2KyiI1qZs54xQ7UNh66u+n4JkCV/KigYUIYUgHhYW04+/CJY7Dcqrs
c/BJTnNefV/eaXGPhi6aVAVYUZdTUQ7t4mgHwgHEFk+mrUs66XQ9zuCZunXMB5cgsSoV/TV5fkIv
EorZe82mMFeqYel8a/vkT1An/n7aMlobWWC2jdOxn4RIaxm3M3b1m9q3at0E02TDxl+AQ4mfPnM0
pVxaM/yFHzBXjf/xpQdP8ENUE3cWfoGZu5kbYGrZuduUp2iCD0am7Amsj2J1384mHPuadz+wRKIB
zUT/KJhhsjc+f1NFlzQGlHCMkbUvaG6eXk0Vt7TDxgCiIlzToDijxC/vNcNnU9/OMZYXmG7k9YKy
t9KC6Ngu70p8HXB/qRvV1gF3h2KHMK+hdcIDD8bUxusbGCLa3AoPHYjzSH2pKfoGxFbWZIvocw+B
58WTXgkxFVM4Ezqjjd6rpbnCtSkkU/LbH2B0EYv/tFp28M8if0pGsCa5V8BFRwVPV58riQoH9Fo0
vU2ck273/R2n11Qmk7T5y/dlgCWr/BZ9Sy9W2SAy8hyEK3V7gSKYdfkGPAkYjSqDLctL1dF/02Y6
YZGFTFNHD6fyxnt7mBD+VDyL73Z8/KnvgK05+qGnDnId4zkqNMllEcPNHquSrNdxp76P7KWuhx/+
9/MYPyJdHjVmnCySC9kQ6NbjhBiLDd5NYa/J6AvL+LKzC68boduTNUQkzOcdtYjr624lRKhVNpcS
Y3rMnga2DdABO+5CFKTcx8Zb16d2N5ZxV8BJjOIDR5/0C6Ip3g2nZC0Y3H1b8GbtuXa2JeQMDFDb
Ye1iFwp7p6pr9m7axg1uXQZSm5M1SJcEgws71UH+e6diXd4yH8d/eSA3I+ufi3go5A9w+CVxgXdX
YjKwtqU5XTp4Plg7fbp6a5eDFL9+kElvohKM9hr0ZuT0hYVP30G0cHhfo5FtniBCtm2gFTHfbJ2M
4xSLxQZvgGfbsRBItOOoXkVAOMYZbBasq6Nv7TEvSAt1j81+j4kaAuAHy5SvzNIS4LUGQgKMoNOO
A/cvz7HJSuGgmo4WFKuhx4f+qFSs6KX5KcIO5331TJKpUAJJ4KErbvT0pfTNVzV8vckiYU1b//kw
n9uyJJmhADuAW7/F798kDI6YWjE2llVB4aAzCirnVIjTyG001lUsdq1ng2FUCe2W4LZ7phNWDbhs
/Z9dj2UZGq0k0+T9RpeC5Y5HHXF7Q6BO//NrMmjVYOjG6PsAhwXsj+VLQhEXGsur7GEMfz9FcRbM
3fDZT+hlQ0fK8n+t4gzBOvGQYVarg8BmrPjZ8lKIZDkXtP5gtIlR14ywgbEi6v7IZAh656mA5clY
wz51U7cKgAUnbXAThanLncOw32SpyAFTqweRshCtNSP898lYidNK4Rqwzj/RKyjJNt1whqn9hQfP
P02ZQuqf6kO5bEd6blaHv+amRZ9yLrEcbgqYPtBDN0qVKZ+8S9suoiJqjp6whvripMdaDpwFuL6J
adkPXaesNwodpcn9RA3BUpJGOM2AhleQFmh29RPTBegHByJMroe+CchXwI+ZanQTwwxCQIllhfTC
FwxCl7F63FlLG3GB3uAXcmFKBcLxw8AaucwAViydOaouvsIsebnoGPH10pqeI1Sk0xah86vOpycI
6kKfayeO1ASyWiz0cwpUJspKLT+durhc2t5ikxsttncr2tzTd5s2ZZP7mrExP0wCnhxdXXmjgfWi
zbfEiWQYQQbXwIm3dekob76dsslm5jOSAeqJKhESlNUdUlCR6LPJJVqv1xfH7+Y/EHfgmCepqvsl
aoOnN7PE5AswJQkV//1yTAC3379EKlsmTqq2ESV0yFuSFK1MiJcne32+hDTiES6sLtym/6Mi3vBY
Hu3ZvbjPHLAW4B9UzumOQ9vTHVoF7NY4Fs6c2/3MP+y2XRkQgLbheqash7dxdAbRlCoh7x8Ep7jN
XPYJqPiIpCH0daAArzJw3GQMc7duOW5s8P84gKzpsk6Zc6sGPUlClWt9lsBs6GwSerTSiuaWJOfe
6DOb2kr5bCyUzueVgOaiBihJTPjqgEpD/20+gruFTonxJSoLaLSP68PHCjHoXUKex3Ink8fg87W+
QEma/2X94OqkvOMHDk1EB+688FS97zHByB1YI/qo0lTBB6F1kty6bAeNdfZz3FV7WTLu48FdGNr9
f4QNHbnwfK7NJNXLLNwG7TF2vyZpiAGk1hb5ze76voBihYDDqg5GY/kWjegPMcj2LNk5Gbyie6KN
x8vQ3QlIMEmpCGg0Iz/oaFQmaxC40kHVDSfzJPmep4hL7zhQTyCz106Cj2hKVonjLuuCxhp94Bi+
mAyK+KO78VhkAFUV0JLAV2zQa8g74HhPVr4BZrW+3OTBOw77zO8JVE3VkAX/VhLJCvyyyOp9+0js
vChatr7EcWyoQa3vl+r2vAaXOK+juWy3oLa8ckGUh5QVcbrrXPSW0LegAfDVBrSphcmhKrZh48xq
w18MwrAVfXDTvHzuAYCYzKMC+AAWhXMlK+bjuxvW0LWLQ7mgxJCWlKHLZfiwejT0ADy/NttmUMGn
nXrrljg/Vsm5OXYXCbBV7jAWKATdpXFw1iE5FWD2TD5f+4Q+sgcEprB5tK1e7BMeaNT76mWwlSnB
hZ07jpYsKMrOgWwWNzlHWlEOMwE3F79ibTdjMy8zrKh4m+o0qPk3TREwMmpGu0+K6sOyNkm35zYw
3f5V43JTkbewE4t5pV8LvPTpPDYs8g+jNU8CU+uco+QHmUTSe9R0zrMtQSJubQQht5+ruEuobZuX
lK378vQnuU7jRzr2QfOJGJU6hLRnxUfrfhdF4VSd5BWJw0VxXrmhaGTJPGVMmoHsFV+QyQsux7/j
Ox4XJqBaXRu/bqSnnA3nJ23uFrBXMxoEScnxjXk7sXvpq8A73FILBo6CJN1Jru1Gu/7CtP4UK5BC
BqRQYEYP2pG0zoWFjN+nV/y30xCXJm32LPMRuqrESXrCHJ9lHan21U9Grc6EJ3Euuj/sZiPLQBOR
l8TwoAajGgbvN4tnT6lFoHthiusJ15z1Uy8i4K4v02KW8SG6MQrr0a+BRVyYUzo85ij9axQItq3z
VfEOMUlRh/eWd9C1yRQcpk1U49viHjR5Wj4TO4hmxELtHch1jfWZC/DbLjyBXQpiikjQToYc0mV5
b+Oo7gv2LexQDFx2252S0jDg4vm1OmwCIArfarCUinUxDejZ8AxiFsCFVohZLqwKDGw2+2x73Xna
OQJqAS4xaT7ezyYtKxjbN9WSvhRmUv7rsyAQIBxFJsatb6eAbXYA1mrq8w0Uvw+P7BInSW2k0OyR
iRvMc+XoAfZyC7Iirl9XvJk6+1ZKYypPi8xTmxA7SPZxLnzB554d673wzG25mz5FSLhkZCEs72zd
6f1+NIHnCcmfhEApFZX69y5WARunIVNPLccjFrFqd4G2b3VlMVDL82FNnwAoCoZv9jTX2HOhQlsE
IDZNGasYxO0CPgDEEehyxRXxrSvp/Xa9j8DKWE/fDpQvFTEbdxrWj1J9uKn0Cj/iha4/6nLyH4Tm
419FsUvPtL63dFcwRt9g9gAidj7faP1CcND8JhWx1QDaamHD0HvnXFMSIBUZ7nB9sc5Ji5zGm4GS
YUHZSTNn1Ah3D5S/F9s9EdJSpcFjTSLIuK4zeRSGlzgw9z87qVVPPxOD9bKLHqN+OmJbtiU/DA3v
UxQVO2gaotT6WAWkyGcd++JBtL+5Dt1bWp8G4dauYm0U3WUiu6SBKVajwvWdxGsfSX8mXrXKCghm
R9TXNticS0Q38YWzumK41TfI6V0jw8I0PTNmOSseYnNjAgBZ4dHGr/OqINTs/sEd+2ijaxkllgid
mQUuzSDT3qaK62ztQ69w35SHLEoa2PbBEn0kjQxC+AigSVb2tiEVDI5rBfxRMyxfJ64ofFhXOLtC
xYczjwUltLR6/AjujDhwz1yuugislmnQ666BX1X2NI/XxiBnaoKVBALUtJBdHOzN98D3TZSWRcs5
NtUQrOk/dbGKRnCYqzlJdXKo1sTM/ytTHhWVIvGfSGkG5OowkLgsStD+GDvoK70lIms/bDiz4USZ
E4/BsHsCC+djc35NCnJ4Qct8wClIyKQRnKTCsBrQt2MBHsNEmJUiTwCiIOE3Oxy418VEdHixkmD5
24CiqkVt2PItDa1iRiju+x4hOL3/RjTGaf2mZwv7zfqhZannyHxu21Fsz+HwGGN5XAfq711+1dsR
mCUFUDr7T8FOx3GrDZFf1rjwhVyJdNv+aoiV33AWjMs5HHjMUyMQ06yActj+N9fZ0AeXBVVqw69k
V4G1enaGnD5Xf0b/LD1VDl6NlDuRsQ/LYTRyK/LtBou8E//8FM0WvRaTc/zHBIpqap/W6aRYW0eF
2D9PfCsoN2rcXZqwqwAphonjwXoCU1iQRxHsZZO2VDBg/1Ssy3BtEYajv5v8hWKdEIynk8CmQPDs
y45ahFomnm0tR2w+1/0H/JzOPovdzg+kLPc/BecRzl/BKU2F3mzAmdqvTdYozB3bg0yjt5a3XJHH
FDSlYEKW7z0HGp9CtcGYtGUtEGOLUi/LtqtnWZpay7FG/bYkcxlbqjKygV2bMqssSXfAdCZ9EA9w
RBwvl944ycWa43VBx0uJhAKPjp1Q4Hhq3qRUhQXOUzGYlHm+zwtb7UfBO5BCoSMjp28XoKi6mywp
5hPdEpCMZO2Rxae+bwtc8uQKcr9UK6/bofCpk7ZSK/N3mzDZHSuGV1Af791fJpvusvBzCWLcL+dL
oBai76MXVZjVYINJECxFcLz6zU7Ehb5E8RxciRWh8ObDkzA5PlIvEkkwnMR09DSs/wh0vmnSxgnl
i1HGh4JKYxLpmm97UtdKV/fHsyL8JyAZ9OnysODLC3LttfMyVHwA0PhBIU7fTrhVnUhnw2aRoleq
jbrGNTW6cfjrteCth6g9ku06R7dHGUUty/FH5WDRKBJq1isxACpsj5L8P3ETBHbdpkIfg6Z+A8xO
Rl3V2YryqiR4rgThjm7py0Uw3DUFsIb/aGnYj8VAoiQGzUmFMfJRZRlStTL/4wvwAavdIsGaCu7L
Rf/LdY3wlJ0KIslRS9ighzojxxBBViCBXS+BvqTC44XzT4CcVjofXaOuPVyEPnPtxXwqL6S9oyzb
EhickUsS6WKJqdc/QKSNTX18ywy7i/yYpcOAxIYZUDQTOx83UjGHvgkDgYKofQSLOkEY41drFT0u
1rCCl29JjMKaSLPylJhzKNGoPGu2d3lzyUVmH8OTmW6x1ZtlbwyEjktLDJ56pROS26bzK8dNp9vE
+eH2cg0RHeFM3+rglkDYwaqwF0XkvKTxcNDFDD+C18cvz5AXiZXTWRa+2a99UZvV3oWV8c0HvM98
G/unBZ/e0Z7/YugKd19uKJGhBnrNcSa/I8rTiV55V5V0Ok/UpndqFaq6fR7QPCE28TR6ud4fKdlr
Hb2uGOXRvd53jHR5/43k9sH2RJ+hcMk6gN8F/OIhZTc6avqXZ7YOYwXMF78wW0Z8+Yud7SrA61l8
xc4ahIQgGYDX7EKMLXOTmMME0hVP8ap0vdeNz5Ut6AZRaMHjdcMiMnnq3XiTYckI+k1VHUP6TzYB
k9wn6Ga6ObVDGs7tEBHyEuEhNBXVx8697GgAjeXo5he422A2kM8t5hALpwDlDwV3GoPzaIGIMubc
BJ4K+t2U3SXSuJTDsQ/lOIfO/eaQ3B1G16h/0kuUDqnxQlXESmItuhFV1Z/XT0uEPFRTS2Cq6h7g
702Xr5Y0Nwn6SrEe8uxmIFjts659xUR4uBZ6Zg8SQC59QnSCtj2PN9xk888gSUr6Bi8Zj164okxG
ICppZ2b1L9lLVvO4nymRGQOBov5sd1/BMcrOlcyMWGLUJ16XoIBqEYUkkt5xho0xcvuZpirb/cAg
lJ7+87mNRjcotThABkvF7HlOFiAOrNduTv1YmAwL/GYAV9PR2RqVN1He2dLFtFb3u7kGH8fbMed8
/jXk2JxNiA2tWWqb3lEIBzVI9mtGal/60rBYRWFws7MjpmvCno2OWVqdgTReZpKtTUg6W/X51b7b
j6ba/oVIudivvmfrdtw7tqZiz1pSF6WKhIQGeGOgYlai3T4qOj4j6+f/0wreSgl/CLxacSDIlxbw
pCN7yWOIgiqrLXWZO4cKgflvv6cF/s+R9duqg18pFxpCFxvY/+CUSKMcKZUuu5g+UXy5uvxz38NH
lSgoqhC7PBVYIpsJ8Oia9MnNw8xTMiQENLQfCoP4GAvTk3ngUl2pioLjlD2GsZvISyNWcIEvJh6D
r4xzZR4bdhiQbl5fsCNYJWMYWkE/sMZKP31bvkVKSe0ULYgKOuGWQaz7RTHF0X8r2D/E4DD2KGtr
nbQgG9UHsZ/1bBGKwZnwXq+DJe0s3cZpaOorQLAQRt6HP0FjyE3qI6sR0sKuZhVhuXkpX/mUMT2X
8tyXwz3ejsKiibnwN12T9iM/cNapKKskEmv+RFPZtwGLpOkzG72OT8AGt66SlpxAv8xOzkp+uFBR
NPudGkyOYGCubk3plq5XDZt2G/VS8wUsvHHtkkylPuvFJNSrewRZ3G1hkJbh9eVSq5eB/RByU3/s
Ij2NmJGKGZPhPTKiiCqxb8aveVPq0cqVB2yYdLFZsqJUy0WasrrXtALd90B1SoUatwd/pubSA2VY
zEuMuyDXlEFELXR+Hk8eK5JkS4/7hYSLiMb6hPlOdHuVjrO9Z9NXTOlfRt6Cwj+zoR9MASy2wWdA
qe2APjO3sUsjo0QeNRIQusqkX/ffpecHzY/dbXV0XuOIhrb3lKhl6fdreUH9fMBJSfBavzzJmVgs
1wz9kLq+qLWGaaf4zLafySCcXAy40dXsjfEkjSKzBH+twEyri//V4XODv0rnmrgHLeAp8jIR/q5S
FfNLIEgZlNdXNfB8H5t/k2L7+IBsbMKosIjhzDl0FG23xD4Lf/wV7F+KBM05qzL9cpc9KrOulcC5
n0apiw1J+7Zf+OPCrEwPIvWp1UXI1hgVvvEIhtlEBKIhq1uVcoUq+dfvJ3tCZ5sf2m0QxiwAKpZy
KhMVGYLZXJqfClWunoNH3RJGfw9TZrpgM3abeuD5pukIzHmE/7gE5jufhEvu0/SeI9qxPasIaUY3
n8jHGd/1CJ9Wt8fIErH1ODlnwoXN+LmmP72z77M19zx+EPomKLWd8nMX96WP0SSKE9Q/zB/8miOg
N0yN0Gtq97kDAJtUqtSCEAxUoj7xUJM2z++K1xbBfHNcXI8kDt6Y8xJVCQSEeJbW7uaaeXC0HPSA
EkCppFsK6COH01bS+u8vZqdd6s2CToRvQ5HBvaa23DzGMK31MB3GaQXg8PBGAvj0zffu8CdWBoOI
AORlH5XTnnaaTfrL5qHf/42hg1Wf4QTNZM4GHEbM7+ObrJdhBKeMn4Zo5ZkaBmD8ipEap0aJHA44
G4vIyztpI8Qdn09jrLrwkpzKj0xWo44Bf0Vw/pnOm6HLOkz0ejr0zDX4aOQGLZMZed3PYHyeaHBT
Fx3kuwc4ubvK3Bq2AOUPWLHrVkmykP5PcwOagkS864i1CXgGglFoytW+yk6fIaQ8PpNUhng1/670
jgfDWQafiZWVupqpsPWL9nee/qANKCB5ifKUrqSBz6DGBhQQBMY1DmOirzBK3tqPi9YSvVpFtFR3
OJ9UBqA6cB/j7uoz3RN9b26TQlYrFLG2Gb5tf9VOc2OWuHfCthPIVqcSXAjyORm+OzYRuTu/SZCI
CuDV/TWPXP7CGOU1RW5uSK7nEt6Xds5+BGiaUbMEP/EIlXd5YkuU/ZlH7sXMTZWeNOIEedgE4JHU
xdPxEVFj0x7TKbuA1u1SL7bE34Om2ixQmiVvm+UM5aOnfYHLZnhOj+T7V5LBHG9OxnN9BH1wUPTc
WO1VoHQJqZq9/HHKYd8do/5K+R8uwG/l5V6VIyTOxy6GzWtBE8kZnbjjElEIKqhm3MBsHIcPa+pf
fosFf2jycK3v7jm8tkZxq6nQCmjCtK5eAPAgIn0YjUAyFSHxx6h/h0cIqgskcLohE77OmW5eKUpb
QxfUry6cHxLNmGJFyBL3H1pn6MwapfLiZhHjiyS+lZmnC25EO6WrhLiaMjb0z5JO9G+XnKR68zdt
pE1bGQYC6pU0McYP/5aaBdo5OYoWiFdYt629mI7oi0coK4Ub7z99ATg8wf2rVNE7BaZLnCaOYUiw
I5cn8U5GaDqXa7fnMRX/XPAB4zDTXuELQ2CSyh4DCVRaVsRfRRkyhndCGZni8NqV9nlLh65wLE0a
vvdK9ir1GsUU+yfSa/V0eXJrKF78JOFDGN34oOzLu+T/XND8eILzLoYvtiEurwqqlQ4z1QIaNfZc
cpMNclqqZzuVwGOsonAqfZt76Z8ejLaUEZhPQsPNX6BfS+LtbRU1ARvYXPu3/M4pAUeeUEMatr2D
rC+wms6W7OuO1g/POKlvfQDDiGPOoN+mJNUGX2ADZqxg8/jrnph3qtCGi6K1BfmCoOLD2a3HVo24
E4ex2Pahjks+nne9HXCd3iaK33kWfsg3bpuVjJtCm+YP6ukZQcjbCAJHraVKeneQhhSBfFOnfVI8
EkPV6+4sK+BlVneGHKuOULSSHRx6SJvmjj0S96dT3ghgLe5vKOo4i+BAruCFBtFT7DtvYFcx8zqZ
afyysw0TWvXPlc+S0BGPqVHrlaNcTRIO3rqOM9vTW813qJromD6r3qtnvAZdTbZUEpRlq1lzr162
Zk6flWak7rX76pf6rtFjypf8XKvTvyEj6/078X5tvqwRNADa1gJbqY6lsDehWdiKrtEb0oL9cO2m
Cuj/FyQTVtM/xImgfEoVkgParEAcjxg3f1HxnvzABSpT1S3ETb36myUulSr0JjtoOl6+YJSeEKjI
1YnNAR5kiRaQdOvHQOkfx/0RN9r9aVkVYVd6snwC1uwZdIF47PD1SKoLc274kLw28ThLuuDyAR2w
JajMmSsb7X8ss3NxjfhLXV5RfFl5gkencWALTKCEEK2fFLbNYgaYCHVjJhRDCPmLpneSR6SKcJUK
Dtqo4REQhpIoptU7nP0yNCNqoKbQ+ATyf2R0Q9U8Gm8EdQ/LTNuvr4i/71TSuwMK7KoubXa3iez0
ASgVo15xluOvepEp9J3evtFKgJzf7Z62+6XSdaGC99Iv7cGT8/NSFT0hvUWAg29wQayhX3l8m5e7
opfXOLcTzwm770zrCXHswHnhiaCR5uRzbYVYl/LhZTYIXsMto3w5mv6NJiP8zcDebWEe+hRR6SE0
Spg66d8mMcEicigY22gGgETpaavjrTpW4TeBF3mQkI4HloFmSaiNCr8oOiWAIYI6dOD+nmiEVPjD
+gqT2i0tdrYHmFFfeLy0LwMfwZGXQGjRWHCOtBvCPRwnoK5hRvCV/TVH8K3H6ffYzkS7dMnAYngC
v2Y2J6NVqNCxAQZLPqNCW2XVXiZL9hzGe0ydzhG4yD8XJrGcCxhfslVpgtMK6lBuxdC/LIo9hVGV
sCsnuKO/lLW7lVAsGw2ntHN/dBogHWSr9Re3N7oZw4xp7u6MDbLq/oqUok1eJlHNgPLYzRXwc+pD
T4q/eyQw5SsPUe5y2hEtR+VwVtGOYkPJxLHuef+OAHwkc9KHpYF4d6dqwWkHXg79ZG9hnWGLmTII
KwIjuCIcOxeKPwqiaI4ZklhXthA3/LdW6EFqaoj7wXq8YNclWWDHd4HFqvlAia1W/yQx2bBo3xM9
+AQBpLp2gsWepBRPUuyv6KefCNDZvoOPCvWhTuaE4kbkjDm1uNJIZ8m9rccjMJiO/lGKTc9rILkY
og6YuydyIpTfyhawlkACCQEmsg+1TpsTPte1BjRKhOcWoNuVryWrD62dWYzsPtQqkkCxhFwtJNqB
Dq/ORPc/ByXyEw0K3TQi3zYvRZEZZ/C6mtfPWA3nuWQkPDOoMgcuyYgH+dSLt/7GD9ckQ+vjmjii
XakjHKRlS8gnmTdT6nFRWpyM3YMy5AYYfsvFwa3OIWLYYbFVVLSoE3xNxIDpoypW0ftS75zHO4OR
d8T3THBnvP1lOBIHCrmAzBbalghRb3zKdf3Y+rcbYEo4MLtDbWTdhnQuXvi487ErBz7ciSjbtNh5
ILrgAXnN0nMbcDVXYEq4cCTqCpdM/86C9qigr3kI8WNB6795hybNqAiVPJgAnuY3J1zjvMqPbVTX
cDl2f2ij5jYWjajUUycAtvE1//bCTCMZRQ6ivmzUwbooPSUKdgVhi0xiWtNWZ/HJe07zcsHpJfT3
mNHZWncsxYKzCd2Xhi0xN7UWOxTBKPR8c4CCwLydv/YOhJDuQMTCjFLGzF7WnuFGdlGK0R3XIZgR
F5GTeO8HoZQ0+mwNdSQ9TDzJm8NyjQ5oJsTMRAG7mnz79peiS2kK0XNOhMTIMe1yZmCoOgML94wg
8TIzOpIlJW/38H5lZhhLStQBIsVzPo+c/bq6zvPqmFzkXC/6CULwzel7ancoz9bicmSiQvq+sNTE
QVHJPoOlADrF9xdLbr03ScPTZi/0wSelTq6aVQtvuznj038Ns3AyCuNw/GM5n/nk4Ggrqz+Qe4Au
Ya73O/onKMsULutwoq1+8/EF6H+O6+6nBknbTlzhIY7H0ccdNTwQMzsdsbirHR+s+F4RHti/yLWa
EGrRH7H9BI8Z5vXlplmD8hB5OCp6fGmg1LFkhce+vfPCUf8mEmFj/IjncSS9L0XVeg5fhROwRJcM
yARf3oVkg8odb2qhJ066MDLycQr5NJ1giQ7UnjdlUnKFjA8D8FJnFVk5905Ob0AYdJhnk6HrXRTR
rurBndxoFC5HdHqlLDtNWw9XDHW4OBN6LyhNoxbyHCa93Xus+Mhh1jPq7D9FMjt7KGWKRemqUHLD
MFVnyv4MmokpfiBuTCfNwt30U6HQ9TEBf9vER2l4gPGPcnpp37KxBCK0ZdbnnMJJVObmbPPzL8TC
A9CfJHk3zBfrg8hKUCIEJHfY4qUc8ByejNYRxaXtjx22zRE0mW0j68vtFX9dIjbJ+NelQJugyc6P
xDxn5BaBsihNa8Q9zgmskv+NBM81QEkpVQy7tHOyDn6zWpESt8qQoYzOA6ulavl+2kix68+0oX3U
pYbdBZfsZApMMOdlOnkS+o5Gn9uHm9semXkri4SCBPmCGKH0pPniOUt1PG7lzAPFklqJIl7ngHXn
fzpmCwvqkQFB+WEQVM7dSsnhwGy2f5hRjbC5xFdn8CmW8Z1JnKs8iw+5TN8dGusbOa3UPHGNEPKv
Gg0CoeLg1e532kVcKEGyquAClR03s4VkaH+TZlxX+q5P7V6h4ArmOKwikAA/UwPMKtG6esH241uR
WY8CibLQ/azHMjB78+17BtaP5dYVjf88+u4J/vdnZixyvzNDpst165Ga5Pw4C29ECUeA9XXUsjn5
+KKVay7a+7ZOIgQBMKINqAOXcDomOsXI4ZYh2akciewpdpeYuSILT/Spf+PBmKmHY9SKxoRe2brz
bb+4Wl3mFBI6Yhw3PjPSlGdT35c9wu2/QT8ZtEOn9/3+gAHnIGyo/degByLKuPV3JBsoMIruky05
pARmelwsuTtXk9teX01kAi9YD2WI6XhiDgr0cOO9e91WpYTeAOYYc0SrMTe6rRq4x8bGsLPHoEeN
87bHn86vQTA32tz9TqEzoZrSYvI57CeQloAau1QEszrMWh1n0Xkylcgnwyx+8XjxX1cwMSTClhLu
JMsMC5654fJTXw4Kh5kO1EnT7OKWe2m62FOcfoJ9IZkdhwHoBB7j8qpnIhMSt96rTpeV9yVBP3ek
iD3onn3CoshRSbyIkbQqJ5KqWWcgFePE8wU4hkI+NuKnkaCQAiA+FR2OmQiMrhTbw5OCfMm0XWfO
2BnubdZXgp8iEkc49wsbMBkfPsejU5riTi8mCC9qWy8j7HQg1lOPr7Y7PTsAHZFtpkHTCMN4srbc
f8f7HftQlwU3Bt0RsW0IQ1WCdL68GeJ2VPMwYGp71FnKcT74VBZIg6+kfjkjOqGskU6H1+7HF5Ey
ybqqbfDEPwMdRrHmmpeJJQf5z2XaI1KHAv6F9veT3fj/hb6O+PfRvoq7gb8bwml5RX8ODm8NP8T+
rIcc9KETPk+ZEurzbtcKmMrCbvJh/Ml5qNyAcn3gFQDCZZstqtFzWciVahIquzPZp1o4R8B6uM4t
V43gEh6vOxzIJg7bwUEhlGlP5dmoTRq2wxPqR+W4SvJWO5B622Xrgg7F60Wk6LnAF/zINbUEOFjT
/ScnZ/xuBRmtf6A1pGSAZTvPPzsW7C0dMiGs1D/BRqQdAPOjBjs9XZv5s4bNsGyawzlt1U++52GH
HmiISmSEr4yxMqCYUm0Xn8eKY/XDX3umXPTR9mj2N8XzLH2CXe64jPtuqESklCTaJQyQz45eUgk9
zX/dKEqZZFka9ZeIRc+8Dicy4iDZraIjSCoIhyziRxCqLKvzIsikxxtl8y9hHsQZa9mERs1yOmFf
TyEnRd3K+essfjnnTpoq0xMKcpi+cYg0mHbIQ3f8XHmtfRwRS8JJikBjzweuqkQYB8TzBoIzFmiQ
NfwXVxBstgQySlpj0Jl77aoFT2zrUJYIHDZbhlGxVNhWR9p5VSMcWv/diGZl8OlkNRVQ9kQTWj1z
wb+O/SjIqVgAM6+DEZPZpnXNHZ+dVlUy9FzEXFUk3K1nw3egKq5tJhbFWrAnTlKwjtVMt+uwWPmZ
L8Muzl+pY4Hmgi2y2JA24EMVQYFXtMRZv5WvFVoRnc7rredcaACBjV1sLxMprWXsb/ff3Ktz3Dg8
QLKhWECDMV3P5aXnakeQX6Ls+Ub4QLkfHKv1eciQn82w4CN9LDvJmFH1FE1F30jGIZkQzKcGd/Y3
WyTLYJebmIOzVJNZ+TQDsRtpkRgQ1RVWTfLtM1E0JaKP8cG8IxJbnHw/ucZ8waBdSYkSUtLMd7Cj
GRxNGlrVD+neiUnU8NmTd3JE4+T05HFJEry8nvh++J/JxMF56ypnCh3VprLO8r/26Av4D1HOxowZ
kGD8TTu9OVDOG3VKK9dTDuCWCi9kBkUIRfA5nEdcK6UfHDYwbBbKoEw6rF2KXFQDZdQVcTySr6Wr
mk/WsfDzaQFXn1u4wbBXF7J9t0TvZGj6fa1xJWDS1c24NinNEPa/OMkvR0zcG5vLYd7TUSXc2igw
6CMOglVmJsUyxmJ3ZRii/JqnTKpUcTZMitxjGP0X0FHtbz36//9ChlgY5vYCVyjzdQPQtQa44aRn
edudHlpE+/GF4Grk4Dnwl88Z31i38TyS6aApFF2te7CbbPV53oiG+Dnpu27ef6/Hop+n9wQHui20
gZCS9OcR1tZCjcqOjZRgpVnO3XZp95UFJHZBroXGBfbhV26E1A3Byd2mhaDReCPSrmn5E5HgdfV/
BLy8rsiHo0ZqGdtUvqF/QIiw5gobLzNLfwab6Tmvx3rD8d/M8ZhfmPQ88WlRt8chRaIUVtjRuI/j
6Ljsw/EsO9Om5Dn/AL7KBHm00oMq0KPEWB9NIHc+5KiPRy3PM2uEu6CcPPgq8HXZZLURnQlsdx6+
tnN8F4y8/QSDrrE3dkytwyB99lxPT8EsW2yfZWl7+XR/9E7SYZsOx45mCMlY5F7WsXzTtDhDbr+n
NFH0pogyesIcZzxOf+hYtCSfyMGQk3fUa4nMnelmwq2ZNEM459YdIbfN9x0tlU1WE1c7zkt7dOPt
Wut1CfVJMPNHWLfKOBdzSLEOJvlGQCswQM6zwhpNdxgTytxVFgzu63vMABdDogXgX/U6e04V+eRu
lcgtdCRwHfXrc1GBlFDV5MdTthvWSO/Uo70lKDHdoHU0s5Xa34X4jbDeVgDPylgYvm3ua0ruNmxW
TaM7q0zbhG8TFyHKQ4bJw6XClRny19nsgFwycEOKjS3pWbgPGy1RC1fE+NYm/qC/p64owlrstU5d
3byv992viUvjm0TK40o7Bx9iz4E/hp2+NvFl5BizPUWXVFfEezvkt7fMxnzw/8vVMf+Kux4B6v6F
v5iCdhOIFRDpWQiyRp8tPNo9wJKvtlDZYxkeMeqdZa5jdlmW3tVV00vN9rInMt+yyxcGJorsrbYw
VwpcfNK3rSmsxa02Gw5hMrRLZsglcAto54GVzpAUHHROHBzxL+d2rNWbFSAhFqRz+h/c8EY7qPh9
yml8FzU/mowob1pstY/x8cyp63P6W115LI4fsR4imR8588EjpSRiWKc8dNyTAb4WUjiD/Qccyn6n
slzmaKVh/U2fG9AmJbR+Dy10sO3+o51bAj/aDkYrjEnsXvfWuYogBQufQjVbBpxq1shz3XUZvQ7p
sRK7L6ky+eTshMr7rE+2ea0mfsDPSmKE4ZXVDE/yrmqCE8scC7IV1O4h4+Qhs+U3e8zYLpVzv8pQ
DgFPjYNs/E/wOQpUe3qYMMZTOJAiX+k6raRUnxzLgUud9HQbcfQ5J3IzjmyCQ7iaDkKzRaIh8ake
q4T+dMyjFZgDwlSRgkBRJniyrQU6aEvR1Lf0QES++rln47eAx/oCMglbpIuWgfjFKTO+rAwxItmW
CHiqbb/XPuKyCT3dBE9KtEwuej8mg1aLZvigmi0/22bMFcoL+FZVRz8wMPU3ZU335lv3VUN587Df
nkSc74cZvQ6szl64rnnIUGoBiJ2sR5hn5uzpD5g7ti5hh5xKVdtU07qpVB2SNilmRdm3T00gwWvT
FQzyVV71H06vuFXjHrVy6NSpDDgmwIjy+cyhjd+l7H5JvPwHMojtjuMhjymmgj1UtbTmSEswEYLh
ZEcZrGDnSZk9WOveNjqYIYcDAGgB6MkqCkC6oI7zBtX/uJl9DtGXjSJoH2KlwHmGc8GmHNq2md/h
SR1a9ty6LVvWIcW6RN+KhGqQ72pa65d2n9J2iKGlPYzD5l85FEwDOMp0Hd4sGDZNNjTz7vOO5Z0n
y2s/89LpWOP+ihXn795xO68q/O3GE4tTRjDUVns2+z+V/X9lPzl9T8ovNOih/S7ljpX7qToYhVyS
isE42AuotkIndFD6zb/wiUwVKPNL6GLJ2L+nyS00z7F45FyYdhq4Lbh8WwTlEcdcELCxruMaZQtW
UwWMluNEbtYKj4TSAT2PxaqzAl6ABnAa0U9av8B4Ea2Sba122QJVc2jnmIHUZUCL+uQZV+zj8HaG
qKtylJP06REcjxHpHmvNqRM+WxCCNu/dCpml/O4q0T9vne10JNOLLCwSPNj+bFQspv4hLighLMth
jGwz8rb60pF/8kGwhdRuABLSuTeOa1++3Wm12ddf1LxXoajxJEtXF0/gRZeZMdsnYkSmxOsSdTKB
rgXS8YSHTrKBkbPGSjlQrQM172BwXjr+MNMPrzcDcfnN0dsJiXirdTKCd5wz+yIeISSD2l50J9l3
Lo7S6kXFX7ieXAAusEYmS39ez/SjzY7wfEciAdi4TUx7sJELfNRShDeuRSIf/K01zrfCPGfnyFhR
H/z4Y/fdeYuLSYORrVF/NrqiE8kJulxIylBPBcv21J9r1IWKULbdPkf6tHkGTPNhM63BqiLHGdGl
iHsmegJSIO9h3kKkzOHL3L5/ktM5hf39TqSowCWQRg6ARVAunAkXB/7WN6vtPoLK4gb8F1+bPu/Q
ZGtcNlHbeeBLlI0yqic/6XwWVy9RnDa53mcn2NX5GWucfqe5PRsg1k3hzdk5tBVP/9ToBNKsci9h
Xw//EI3pRPWRMB9+aRnJ2RBiiDE+1TyftJH5N+nrN9NaxBCG5z3FWbhAQxb0AfFnvR4T5eX609nr
lFAypNdU7WGWr6j9HLxwfrWumxjI1vMoeWl3daTMXion7CiKvn66VX6G09I+/FRm4lC+CWQBnxP0
72+jzOO9lXf4w64NP27dD9SWZ+Y6Yr56bgzAaH88am5cMeGgM6uywlxkdvcCBmNIWf5U4K/fkxPr
hjAIUrtRZFy0Y6ky7xgIdFIAJcNieUG/bLqTwMiPgjOMLtl+U+/IzO3ort5Dvp5Zm4A/RXc8UIQy
chVqkY2edU+r4YadrbViGRvRWM+AwgTKJK7BiHU9MTK7aDCemh/v93t+vcHTJJ/Qu5tWBzdk98gA
g8RF3NBmuhLaPkHiBv9U290MZKLlMxhk00OseKkhplmhQfnKBRgKJPJeithiz6RMHfFxJ7sMTsL6
/z21WYn/DQPNUKHvQaMlXN0dIa5frVypnZBavw6uJ6U3veAtbNnk5xJ2PhdI6ZnY/yWIOeel0Fhj
EuRhdBlKondinp+1Ac7eqVyi/7BllNYRI6X5lpSOuk7XogFJkJNNla4b/Fqyr6Ce9vD4sn2kMFA4
UFeBemL3vJ4xqfCiWoGzzz8D7VEALkmXWzH41TDi4C4e/3722UVa86V5RVwuE71ot73f/Tr0GLx2
sjh6dblihMtKOT2SrGCA+BnSQZUjJPK5YNWyYrFMtmS2WPGGW/3de8LgBhyDU6nuH8+O/DuYlH/J
iezOn3JzCs6nGfI0Np6KaFOjzL1v0Pm11MhB2ce8B7XM/aYFSDVgSTAnh2qdKbFPGC/zwikUTbAI
H22e6eBoSZ7qCS1oHIaoOlckjPkd19uKwO0/QmWe4OAOy8TUUVsxeiSf4zwQPxm3tKG+bT6TIkAH
Wfj75on43M/e1r6xxTtt5oy5Fk1ZTkdpA38IsCr118NTKUkFI7ZaMsQu6Qy9mF1n6JbQtlyXv1zT
X1ClMXH3aBSqJTkcZhRdCU9yIp1e0F2KeIDUW8HVhkkASyybweNI3JjVjtJq7T5KraLWHxpTDXb4
HjrfZRXoh8O4Wg5T/POZk3nJKH/MeoQFT6N0qOkD36+0UR293vphGsVivinL9Hzmb5o16egh3ipD
UQpdF+LF53QzVQIeRK425uJLirnYe+98OgVCuBFQgXyrPGehdA5VFK+GekIKw5kMWQLyzwaWrJhE
LxNqAWWwij6hckbnYCfzp1mj9qw6t2HpXaleXOL6mBUGoY1BW4tNHnfKJtL4xKbLw/0bJpW/ENhV
i4Sv1QpNd0tl19Mj3G5zNsJvReReGpT5HgfOA8C0phLHqrsQE70r85XctH3UUxbXnf4bYhte96vy
PimFdm4I+Rh9hvcUBwQVDc/B5FCaZD3QfvFvszFUnluk3fbcKNrrEMLWj+OpT114xl+ErycWOGRx
niN1Xg7ecUSoFXwhid6J2BGRahu/THoMCl8v5FWV6VAicCzphPeSCq0OjHqEnqtcqgPrrK9B5bGO
nIggttlYCNjwRgAsuRVuqkJWyD5Q7+cUssKV+ZTr9CTuTtN/RmU7jJLRzhHN9CjQb4/6M0tLYQAE
KtRC6+CyyDowwu6tAymPb4sfpXIjHNWw+8kdLjGeBiM5Xml/Q1FLSAowBHiRU/etht3vNpDtF5Qx
uuq4Xr6rf9jK8QkHBS1Vuas/Xuxo3u1hC/Za77sUTjLT3abDSFWymjuMqaMjaddYl4UYAz3KyR8D
vW6AUC7I8GkwwlIr9bzCcw4/21oN5nMXk4W9tbaMEFknPHy6cLzUJhTmNUVWWTAMmQPdPnI2lfFT
IjhIclsRP3oJ9HAUAMGYXyY2FcPMvQhbEpir9YLVZuYKmnnMOIAEmQ3ACDVylQndUHKPoMaWk7tY
hp3AkkoKzdqcGcyc1ASJVkHdrhJzKNFefU55MJebcmCOlzVS7jZf97D4XuB/M2FQZASigttglluB
j/XmqME1V0fQChm4q9xS2Ms5obmAVpJYRm6Y4Yu8OpqukUrfcTpKcSeYNn0ri2dnne8W0q/zJgyA
0lOpYppm0PbvAYHJTU0Y3oDEC9MMfCo6iuzCEjfQhXy9AZ1siVHrys6fmoLOOg0rl0upEViDzgUD
ysuaw0T7ZT5Y2TbB+0uk0tcH/xlqMVTQF2O352crHByB3yavdHj6xkZwxFVH+uQ/TEeti/fESs2H
BDluNg2SeTUBHhX4ANd6H4lnv2Dv21DmymOrZXcvvyTaT8BxENJvcymUjJFUxOxzR4lUNcFFmjGB
rslq3PEitt0l4uqMKbVnVzODp9/THk9UZ18zIMUxW57nelcQHjX72LXRmXg8btaVRYYs8SLGiR1l
eicLIaoranGisB2Cjg9w5KPLbNFUfNIBYRV1lZmZay6e5VwCYe2ka172saHLGndD2/fhEnA/udJ5
Brulr6hPzMT3oYx8SfvBCiHFR3e3sULxA8Xx/szD9QdWHP7TXJQH/CZGciMH5eCjPiDbJ9nW0blx
Zsv6szQzNzkOOVLkDpXyQAjcIACszmxhrgYzXHys1e7HMJ/rr26eYq1OiHPBCYFQpdYP26xC+LPh
qm3GSrPm2T2SKhKr+QCbw/IDY8aA264TcSaXqxXjDkxwfJ/toCnCzh6g/Ax/qWDA+ifaawI1fenq
v9Trx5aBtfUzMO0QoovszYL/5AuA0kosTv0IpcbC1UyvKWSz8mgDaYJnxWn9HTdAVFlqwc3cSzKB
0EHP10YtEQrQCW7spPbGwZOAmnc4QF3MkceQbBWCRX4MD2x9Hk9/d7NFXjcaDEE4oB+YtgyVi0sj
L0wwXQNhl1A7qVM2887w3tHQBPByORF7TArRtifEirMAmcwDXN+FUp47XKGbbL9T7AQf5gANLxzs
/7Lwd2O8jtMc0phcLrQQt4vHWBdY58wzqY3ZMPL9+ClxnJC4TnOfi43nEmd1cvyDALWRoBs7mXoE
Q2b7/gS1HqlVNZzR1WLGEIMNSU6yRrEgXzZz0jGPrMtnNMeYdAWvuPK4pLBx7PxcYc4YUcoqPba8
Pc30hFpdUIuSWUGly/SJZSJcinLu9yfZ6/GsAn35f9fxvPog34EVv/SJsxJqZjm5WOSRAnhP7Bj9
l/2xTwxtYN1h+MgHHVgArYxfo8E0jURWgceVw6Kg52rn7fUN5w94gUWPfMewVmbDKD2ARwIe7zE2
rJSwzTDP2Wjaooj0vaKcsplucqOu0svQ5kK1F3aHiNwfLmX5f0EITuIxLv8Q1LEoLeFWB5nLPmdC
825Mt6GKBQcvXTePGu/1yDLySyxvPULY1/fOXnNxIAQpb54uV8fyp0whzCiR6JAKa33HlgbPXzQk
KYPghKfCyYkHQ/LiNrvF4jr6fHUjxk2H4KUK+XbOB8wLkJuKYYiiRuGQx9OCX/hhiTzp5L3g8lF+
FvkRvt32oazU5OpRQQADsAE/BrL5XA4iyebxUYEUo/plP6qFDntfACGI7bfll0eUQjcHkGPf6c7p
4Bp6VO8wgbXaM5dSvk/SIsSN1HHeNXHunwDdCyRJiu3VyZiwzZ1lZcw07JrKJYoY5MVII6XNq5DF
kMMxH9ih6cmHwfcnt5NLvJN7WKLNVqo7EMn/8wFYx5u1ne53F+l98SHzFDtbFOrkEEw9Hg+6J5Sf
jaKZWNW1veJish6v2E7EMTCD3a4XiQ8rHr5f9N6ZnQyn9KUD5tCKiy5ebEZo8lNQ/4hsCkQAsfw1
ub5e968+SJyEedC/e3cWW5MSqpLYUmfoWYTnAXqKgcJs5BMLTObuHbzVbPfOS3NE7TGl8ZGe5AiV
r5PuwwL1YEbA/t8l2R2XMisLOjYWwS9tT8gDljyr+rsgDHNnFbT1fWs5NUMzuNnsAAqOOkb8v8Ph
OaogbZJ15W9Ym6W2EctJARgKaMMgtnzIfYEVDwoX+CYpszZgoDpS5ZFqDuMQ35EEyf7yXcteikT0
2vh/PKgdEWmFd0mzBHhZodp2+QcZEqrMpLGGBr6pEtjCj80p4gzkvVGv5KBq8w/UEiNAoLy5aWWE
yLKZwNUuB8Bf/VNMsBwZ4Mlen/C3amD6SfTKgoaZB6NysHCIHl3xO85W+5bIEk+Kuq5Q56fL2O+v
BLadr0oZ4JG283hNHankrvoACqOBTJmmUJxDYeDfYxoQaxF1/gMKDetZszjQYHfC5/cKe+50JRlg
cU8ZiGIWs1jvbluunFLIknWtMj9BmMhtGKgngPb5c+Wxkr53wEqrnTw0qg/CCKWgClGV5LUYsK9Q
I9ubv4MU+nzwGO4L/ip7TQAFApPdDNg/vTxBWqgTueiOMUo9+vLU6YXj2pktiERBso51GhPyV9LC
BKBVGRHo6xN8YY2j+l3pevvYMI5fQqPgxck9EIJp9wmVl4RJN8GHPrEcereIVPuk1XShxqK3SfeN
40JtDES9RwLdcWd0KAyUSR0JDB6cRKuX+7sT4SX8rROtURwddZZs6G6iK6jNeA8aYRtTBSLE4BqM
M1QWHDPb7Y3/e/Wuu/aqaK6qaT9ZonHb992/zgrEGzHNPw0zhxFm3Pn4qU8lmoTFD+1Y0NAiFJTJ
n9pd3x1nPwvdz6LtMmGtDnyDPNIevGVJ88yo/qwf0dgWk6qwGKstPCKm3Pn7Qvv+wq8WZc5pFzBR
m9MpjhdXiHqMirPSQxKVgynH3kfGWLZaZeFhQrT1GH0S/SaTsa2+wTt9P4Bjkn/2Bhcyz2hWKSEb
+0mIlAKC6pxAQKqNNQfcyOblidGqb6KAZLcEeaQycDsCBsjoiIJqLMtERtLR8VMx+um9tVllWLfG
O13q9opPaiVyRSSNUNv4YdqEF1SxJQXOrjvTYuANVQ0rI78NlgRaLfIl0V5tkq3Vbbt+rzOavJZC
9GlSlPOsAkyUKK7hXMEC5Am6ZMRYQuHRPjse3qhOHcUJ5nYlmvQUWy1FnEYilBIKGjZMxq1lSHch
6lhMhMEiIY/0C1ycpsc5o4OXtvRbyql0Mq0NZZHocKHTzFy58vjyuNZvXMz6iCF1ZachSCf/NS2j
Pt7OOT7uZtxTOz06BrzZC5mXBQqQYRC/Q00YaaJdo5S34/gKqgEuA8MSqjjHAfoIyo0mMPB5uo4O
fl20VoCf8Sl9WZWGj8MPzNTOpCnCeDVL8G1PEiZwOp46uZoKmQ6O3CiBdkyoOKH85qpY+kUfHyYu
l+0ynek3bFYTd0XydRBhPUVAtadsPpxzvMuH0fOdW5zv4z+LXLbRaogQ7GftidmTQrFZNK9rNNqB
BRM1z/iIpnWzs9VbEbCBDl1tq7NiMgjnLd2YnPer8e5kWM2xOpZGVryDX/P8PRxfmADhsMOjq6YN
P/665T6ML1oOjzSEuYRnlFlp0AQAIUtay2NGbywgp+lR8dCDIPYVNu/6KdJ9tzUskP1ZiKGYyC0S
iYg/Pk45W5nwAyn0KEdaO+056A/auczI66Qi5JfylIap+0k/ok1sSUiuhXYH7KipGYPc10SCmSGj
wKbhylaz0VSNWsemK62/n8YtpCR3Lsz6nN25Xxlx4eKKwUn9BCN/M/TBRuMuflSzdVUB1vpqKpN8
E41OHiYJQ3NvWKrX9yyXqYyxjiXDPX2n+QM7lwrb/tBXIa1nIc6Fn6ul2At3hJR6TjCEW4OS6dpZ
3RAIOqSouJpCZYLEFjqYI+sv5QmOUa3VCcZH5nk8KaygQ5xLABJ3b9qI0pHZG6VoO287NjQ49YmF
6aiB91eSTLwgPZTqWEv43VMnW3DD66kR4gr120IRwkLTGUY1CmsWvR/45GB0FY+DI5Zf4lvyR8AE
2cVHOmhfcuYfkG0I2Ujo3KmIzVz7tCX5ddTh/qFVZZRHYK4EZ7ikWO+RAt8k9+x00/TK9htFcx/9
EmsKtDEk9o6o8bYq+yJtgqzt7rmQaLsfRtkgsN/2ocniudevHU1+IVVPWLJKkJ5lFiwFbWmQizI1
RXnsXCvWTp/MNQo/y8LNOEtRz4/tBPz39fNkBL5PYf0D/DVGruHK8DtP9ZcErLap5SIK1Ib3s2Mq
UY09hm7yxrWq3af1ZYGiu9HJtHbit9CK7SXm/Aij4h8bxtKp7j5B518gJSmIxT3dTScs8jpzNy8C
XWP9FrytWe1OT0ik8BaAOfsm9B7oJyYm2PQldLFQSlUKLofdManaMVXJZxMr4LYUnQdmnd9gdhik
hcaSDl/jwWpjLkVnqxebCguvIRPhiMjbfJv7FO/wihaPOG0+bOeqMgwl0CJXSalmhu+0SqQwflLb
XVogk4DpU9uGzsydaspdnpb9VjGrSg2BLf2jZjCe0uZamFgrsh23ru5c2I/ffsT6xhfibgwluQaY
Kni6fidlJyP5uJBJ2dXRMb11pn1FCALSXnykAyiKKQMiGrl6LAe7RZNBFJ1xdXl3qvbSD7eYOCqG
0t+W5puL/Z7YxihTCrd4u+O0OkQ6LWkuyhDbIDX+5t6uMLHVsPYE5KDbkQ07EOO1bsB74YqBwqdH
31lnEOlOcBdUJxK8NlwLWsd/AcC3+83/NfpXc2TaB+hv8fxcGI/OWcRRQLMvr7//3ZgyrtGz9bK1
CANKbUlAjCrKQhRG68zIkoZbJAWWNIzgrdk+tlntzkoWFOwsNnjexVF/dJTphCeCyZo6dsu7Whsp
gClLz6cMH0natWJxHCSuj6OmtC9NsI0+s52i8XpJLFwoW0ehSXpAxHVbMegIRhpA/2mWI1Rt4Utr
dAWWLIzzJ2v3xy/nuT3L4loK/MKL8mjHf0qn6tSWAfiaOjJbD+GZrYZVz0nuR6OQheByYxJqMjNd
W42Chgn93gd5VsL58MM0trT8BmFsyQ+0ozjRiavJ8w8gJIqfGF1GDwk+V6FJyNKprdws/DvSg3ig
cKDccLuqC/AkxPDVgfFnkQrM7Jo1qLwbw8LKXv0mmrv/T1/5TajP+VL90V5yQt604BXSKO1utQtj
ZWWVDphVNtd6MdqeM0bZJjE080G+FTqLIthZyJ2/Z9x0wnag6WwZebuUOZpZtyq5KV1vReV1Taew
9/n53YgDvOzEqcKcYaQUXdNO7+jQw0B+tzr2unIUX5nVha6gH7J0oLJWgyCz3a+g/dy9c+GCawOt
xaR6RENXtzM38v2oc8gefFvhxhGbEd9w28EpSLeyD5YiVSLVo//IugO8vddQZl4ggb9JqQdE1T3g
BtOSid0us48s8ayUZgXu6MUvf/9tPBfSziLmkHJfMANddGGBC9pc+FBGVmYCRKM8SgcpNtpweq1j
RW1UZe11/5O6ThzdqTOyibn+/6lknMcvCv77Vjo7lbW1vZLk0JH2hFgyoRomSuGAfLPlDiPEWoSH
c4ZQbPBUPwYIcx2PmA63Jm+VNc8PhKn+Ye3ALjgY5qUE+Ew7V4wQ6EK4TyLYVfnxrnKa8K4O3wx7
BAvQ6AnfjM/9rGp3cywPPt4dWUrmOj5RMNpJyswKRrTw3Iw0s7uE+z+QgrSDu7LThuasnBBXc/VD
xC5MUIlnrglL+qwXiVWS11G3bQkDQWzRmEfgM2AfWgAI3tvSB/1P6PqMIzgtmehrj7O7U93ups6H
53lLRbUH7hS5Voecg0oYH+9swuGH2X88vjvU1tV/Ffpco7sUknuPypNYmuJKlSzBxRASwikxYE3I
4O3/JLTjBLYZugQxJAHMUhOUwYAy/CGK0CfQJyYCvQBTf55yzePymzTKISmB4u52Lcy6HZ4DBrVT
eltW0zetyB309iPX+JwuRNLPO827lx8njVWiKDOCZGtrw3SNHTuGj8Yz6Puqwl4ATdIqau93ne3B
sFD94L9wp31RV4lBwgok1nw8lTff4Du8p9VGLXtaVZbmo2NAEdwRjAIsnQ24o5ZugNj2kfsknQFd
J6lNRNK93UXv66zyD44HC0YAHw9FdvJDLoKHxP91MRBSekPvfb9Z5mE66fPacjusqp+bh0zd761v
ndqMYl5i6CnLUcjHDFTVG8ECCJ558WJq91nRjT57/I4uvCmupSNWTEabLoEbuaqAFSIXlsjTaM6M
sOjhvAsh53hMSQYVSqlKfRWUSZP1+0mg6qeu3iSkMMI6DA1sXfkadN8Zqkqm+ib4YGCyqsbSl2cT
GRkMmwqo0VWb8E2aBpA4Obred3ch1qhJUFGR83QTppDShGKjumV+59pu+PVrk5gPC329lNEL+3K2
lknmXnfaoHPMMLV7CfFh4HNqJfTnvmyclBhi6qYnGmJe9QCgAvIBvOyEZMhHUeGr1+Z6SP1TvPf+
XNJMpgySFdKFjdNDf1YrWnSSsxrJniXtde9SoGJ7/8k7uXQRZjL5d0NHYFeSe6V5U9cge7jaDUeS
lw/Ubh84Mb2ogrcPdt3VICxNQjNCGwuYf2Au20CyMOdigYVtgus8AUEih7aYn5KnZv6NkeMlF1s6
ddHAfm5urbsiZXWtJgul8g0C1+Pfc2TCjoeLaEEOzWBlx0pjVdHByMsATSXZQGoOZblEPwuKbZIL
bErMGYkC6whc4HhHjVbnb9DTa1AulPe71FGIq/IOgNX8SnWThWiCgF7o2Sb3AJMTDsVVxYy2kAow
12WtPF3pmw3BX0jrqUY/HfREzj/CAQQMTygR0ypvDpN6yRSD/BXjK27Vuv7xPbmzuPld2zkw3cOb
a0wHvb8r/XZOoLOMOVvQ7R965aTslKNiYT1EUk+sKowjlE7czNAVzeRMLfRLmsv92XmnEstI71B+
5GiVH8ZNTPSI7GK0vu7E6QG35O/XlZsZqDYmKmfwKPYKceJSZxPaYu36w21ILgwKuzW9p/wdG//1
/uL29kUeWNnRQVqIzcCwkP/Bz56nEP0FbJ6623FlcxNiDjwBQR+kQ2PXjqcY+5QNS/2SiKJbH/Bi
BHOB2udFyPgrtk/v1c/GCMoYORKAAbaZddTYLSXZohlaERTBz2atlzRKWc5k9EtwZ/B7QdCPKLkm
6R968LssvXIGzOWBWwNjvGw0d8FZ/Vc+OpFKeW5KktN4OaOXo6dSx/RqscyykLhlTL3xhgZz6ubM
kP4KJgK5Ot45PXpxreULBKv+XO9HKGJvlLp9HpQ10QGiJxyzJ0nntUnTjVIpdna6R2B+PhoFMOSg
naVNSgZdEs44fB/8QdoJnxQH5ebhtISJaGDjHBYbCnqctKSqVGAVGFpsllRW6Yss946E1/c9cnGd
9fJqgMX6PWs8Q+7OCXFha81pfgjS/qmUDCiosEIbTWbvWWQOSo+iUBXr4o68m/F4h3bRaxSZODMC
Eo1jegTxm90YL7brTlqub8tjBewI4cLZ0uu3FMM7FqoTIxnZekoel6v5OoGWiSj7XyzDZJdSKnRd
rdWFab5DFVU33gfVJnw3HrRbDEyYZ7wz9XDfWhMYj0sHDz4P0NA/0MA914qAfCk3zGU/xoK6q5QG
KIb/XurNoj556PQ1w0BJPmRb/v07NV5V0lD2LDRpbK9sW6eIU3fxIctN51MtSxGJ78MHj3bQKB0g
K7rrLDwpZLlQZnMiPxLB+Z8AaWWmQVOVpG9MrrUsPYEOMC3PO71gGHbsAjkQc9C73dWyy6zONe8V
jl4Q+4RAhD0jRY1Wfwquj0dziYTJc/PKD9F4VR1c26FqFMuGqsdsKOCiDhII5yFRnT7otpoBi253
1nciKRZ/9QyNp36C3iSaXGCv/0GMZoLE0BX5SyF1EaUDII04+5XCIRAew2X3OD/EfrqkMbUhXdd9
69M+OxcDkQHVcj2cEJRRCIqdg7d4yUy1DknGnOAC19aB6jZYdmqH6L3MtpjP85R1xh+dUXPkD4kx
nZR7FCxCi5fMvpLRn41AczLCKNRBRGw/K8iFtXIuy/dYFhDPhGVyfmGKrrbsa0EZpdwTC8Moniu7
iFw/NGDE9b7EsEWQhRPGq5/I/P9SmpBvDbXsf+Kgj4FJoEymsPg+QYsEu6bgDtUYC+Sx3pxT5FYs
4hR5GsEn9xFA93EVBd5W4jS3GNEvypE0k06uVLyFQGQFMActwpyRETOhcarp91+FSGDahAFXdXtC
Kk98XtSV899hKaD4sKBlyZR8GHJVWB0XHFhRK+37FOKuXab8IYzYVwmbd57m76PH3V2wAzL4T7IU
FRw9Wzh7PS1XmO2iB+ozKW4RG4vllsCg2vfHmB5zJ+dcFql7Mj6BI3kdyao0TIwsyy8G6mIwMudA
GZWLAOUS/CIM3fEAwaq9Sgcd7lzlQz5oOIwmYe5AJLxKM5AijpI+UtWlf8sGmvLxzF6kIMsTgdz9
9whkRLmubFTxW5sxTHUaJ2r74ZvOETYhGlH4I/PEg6OwutojeiGKTVy3uUrCWIJD12/r4QX7VB4z
8vv661doWkIpzNOFKp/gIqugz488MDr8jBPZGUs+CY9is7Y7hc/YSmNKDZbYyyw2Alc3PWyZvG/O
5n+18juFq/GQ5FKR47yYuyebc1txVzOy2VKtb/b3kUuZ14NQaRfF/ESOI683sMPrd4iXX3Dk4COA
Z5AzatU+FTjHfhEhf2h6UqN3hd4nrk5qoAn6lxPtIH9RWp0n4dynJ8SLLbz9tB8UMoB2DPlHNzPF
/1phNL9eVcCwDVm0kilmalELuDjRVxY3rB9U94CpT2PqavsqoaQU99ewfp0JrguzR8O8AenfUhwJ
ph7C/qKxemAFau3V/fbTMYJyHVJik0bLaEFlojFo6LaCoGTTmzh2BfKD0vSBWsf9/KEOH/SX3A+b
F5haG6ibjLngdwUp0Y8gNN5jop3t8sTF4b0n5YOIQSxQChfwGa0yxGNiFDIQeMiXnF62ZYloyiiu
7c9eujJL9zsFskcuviu2Jfppq9+hNmJNhQNEUMql+Gkv/z6cKXTEte5YiqGCtI8Puosj+R1Bqaf+
zgHV65VXpidmRjZwAtPFYRTRw2D0aNeysg6e4tLltS/5xzyWFwCRLAQ8x8qWbnXMUKRtlOD6uNW+
hCECIykfs6PaotiN97hIJu0A1p/loJkhstoiJ1s6IxIrQ93fSW1sXMZYeKbPw/hMqkvCUsolyPAR
wVmQxA7UERlYdsDD+pSEGArh+ErTN29C9CtEs/nsuUhofKL0vUIHPP6kSMHdXdhStzVn6EWeBsnw
bEQiOLC2oaInbuKQXLxNHWjIsz803UG7JJ93oTYqQ+2f6Lb/U/WWc4mtnjGg0QgJAdvfOKya/8lR
ALEnIRfIPllTA5sSEB7/PyMPew5UpsTqyEXTP/rzA65Qz8RDJX9wFA7+ouQM2IEUIbPMQzE1pZUz
6VKy87L/4ulqQWdeK0sGZrV8pkPcntbyoOPJFamMCxSaJnYpSTBomZGKE9UEa+A2ZTeMTVkoqk59
n4Gpvd1JPF9lxGTYC8WKNpMR/1YPQA5vwnzHq0JYLT7MHDD+9+2O817Aw/73N1QmEM7uaKPkx+sg
BSRqJbPbZAEtljxkQ+jFulNH7t17BYOie1v+hMWuMGl/LGcZM/iFn/sFgOBGYFFkyPtyAZv64Z6i
TS10YbdH+FE99v06VVhi/rYHN4AUByoXTXV08br5sCNPTrdftVgF/LM9PYHGjLy/+wayvfTcGRPU
kSzcVdXW+UB/TVnGY5OWW6quLxAgzwAmKfR9Dtmvxg6DNchfxl2dXAAZczvgdVLntziNTPqDl1w4
oS7d7VakJaDv3KDYVVHd230PrlE9BtVD8Am0u2UKrg07cPFeiK8J2uuE7/Sol1eZdcG8Npxk/7nQ
IBn/Wj/HauMUusYmuGCS1UHnSa9chkPuh70RDMnMs1XfLzOoyMT8QnSWg3Qw4Z22tikEaXu5Mm7h
/Irge5LU9Ip3z3QevBuK3LausCbFgghwnwXnKJ0dfLEaZduhFqzFzYyX6S1yj16Q0GxHUTe8hjrN
1cHfmHIZOJr+kTwYkZLJPmkhj60y3agDb/WNix2t/IyGTivZdcLV/MzrihMQJgFi+6wyCQ6M1PcU
L1h7KD/1wpUA17MxXaXyUy932lqMns/mUQ57CyQg4qQakC/KARNn/Tjc6OEHY2Un5leQNX4zVgxF
xEqm7jQyWFJJL/IlMPRESdCsTH7AsImiMwZgnprXJZz07Gt2orPruQmNrdfK+3umcYFNGCVhlVnl
ySh+S0sJDS3QY/VREz9q/8owrhJT1kCSegT8y2l5IFtynjcfap6UAw+1wyRC8CKw0Er9dOXrDzih
2bcyVyPfxypp0s6+VhOP2ErEIMTQWhtvxAvUn7+gohIsWaTopk7ByG4jnw/D+f8E/8gmR82vOj9l
9u7OYaTU+oLDKTXHkWqVQGrRkSaHGV2RQDMHXvbkEL6+h3m3oq/Iu9Ns0XhAvEwDpA04gjyiRrGx
JTBi/SU7y5uMLo0Tn53m5UZTCYf+ZmqFio1naZSfI27qoOpJLs6o89NKnxAXAxA158D6V1qFMYTD
1vR4cV7sXIkDzpLk1Eic0iRwiq75dPONS2CpTXTcI7hn2j+B7KaWH3AbJq/4r0UUrnbVQvrFm9n+
xD1D6m4YPzFfRVa+s3evfbrJ6Rv2+68xjQqcAsvUTDOMien0IO922nrJ3A71holQ6w2LOydDuyAV
MZNaW00TsRt779MFT4nTWNCV5u3a+otOrlF25iyTF/+lE1M9pk89+hZXei2okQhSP3E6EelOV0dS
oR+7qOH9HnpL3Tt+NFk33oWfFkSSlZfWg032e+KNyaLuK8/nBy5rUa+4U7JCdLLip6ZKqlD7GSHn
KgYSLcPBR7nicjnP+qTizB7tB7hbQFQDfZOLX8VG7yu5ISEBuHd63TvJuEmQrS+9tzdQypMeSa7a
VfvJWJH821f3uOtgZykg0o+aOGpEQbOp/utxLuY9wCdOFHvdSQ9HvrpXkdZhB+6x4uYLcF5tmCRI
iN9LUA55WemxDjjVHakR0XkSitaYE3LSbPfiwhEgQNWeKeX/2BBGcMhKfEu3spwVzDclAlXJdJgm
mTO38tZ05cIOf1YGUKkyGnRe/dCJ5C1pEn1Dvf7IJBz/3PlZ30yqN//v/MyU6dT9sWBxHfU7q5OM
kB0ZfcKQWZFcxRIsd75O7kNi11N7FMZmvYHzXgARpke0QfTQmIgrO9lMviWLA6ENAVXojgNf8SiJ
UoFRq3dX9nAmjncZeZCRwcSA0m+y67Ndk5wI1k8PPDVPpnAyBFjVGaIq+EDSRpH2Qmb8//nZPCtL
sWO3TGj9Jxz2XVnnYZjxcLQIel1jk+ZTlcjPL2Aiow4TWgXa6w4a6QOPI//0cHgDopSKEs3m1M++
AEPathGNNeNlZZnrP/x4dsmEntsO7Nfob04DWo8GZg+c6AfBHQx3CLlQEkvfCNIjy7RBR4iIV6ik
XEsq1s922h815bvjp/0F/6BJuF29miwfBNt7Oa9wsGqCteRmO8dPP5zheOsZBZQzHl9ytccnVKLr
1hs3xHNkjC+1gsQZDTfjBQuPbuA0I7bU476V22TQqjaudRkLnN1OoVXHxjb6usMDY7f9UCYDjmBQ
tT27DDMhNLMvEcS4p3ei6gSLO2Q71XgpSldT+XHad5Zvt49rjP5hDMtbAoDWij/xxsp8YhmGOKft
U9TPZZL+OoUKALHKEC19+hR/2hAIwo9tF+zcpqw0XjzukRZz3PtwNvIGh7kyAg2nlb4Hzdj2hmAm
duc/kFFR5AwN5mDwLfnclSnG1X3YhnwfJTDEeK7AAPULB4fbiKlqFOAtDOv0BrY8hcjUqvSQBZM+
3qDPsjhf+a4jmuN7gG4Zr+1efmPZ4hHemCWWLWuoezDres7I9riFWsl2TgwGEMJmUmUkyPj2/HEB
blCMaMhiYrwH2ZpcrkXFxs5u7kR7KLyk3yQYNYonnrY44aF9wgytOXsn1T/o6tuZVbU0Z8+3Xwu7
cFBYu1NHzIG63fGe/Ldd4f1d/FN/UTMF9UxsYTiFejE2BsPh6+rl0XzU+Ct3NnGXXHrFQK9tAS/7
EdzIpW5/PTkczukKx7OyJ5M6iPbdkKz7aLQL1hA5OtOZuy2NjiMNaZtoe5mqBO8K0i/m3P916oub
lzAxO4eHasljaGmkdw4xfzn58MAvVzw1JF2ZS5CD4xP36yVwq5skHd7bx2SnZvL1WDpqsAv6M6ri
VHSx4PFcb3PVgPNc+N8sXv5Ig3OSaILntf5g0rcAlTxMo3wR8PWIhEXxjC+/qkGDk9x4fL2dovf/
PBzTv/g1ua0SGgSiMNs2tXNvpJiUCR/+2RIHS4DDtgvERrF7occ9jBkEP5ErIqHELb84bdUf95IO
vMdtfZWxE3lmLwUWDK59oAxF88uHa4AkE6JL/iYe4Iffn6aFhrYp6kMobXd7IHzCCfNcdtieiQ8U
kcli68zNB5bGWO7ovgBvCMsQ4MMUrgFjUD8vi6oLvMXGOtiAZF9+2hjhtnlt0H0cBfWMcaUhCvBa
4WG4hmREFmjyCZzK+gU8aQG7S7Q1c6qRr/lcL3N+bOyzE9QTwDrfHMXSQHi4aIwyMhtkKri9vtY+
m1lPAKaLLkl6qjw6QeelA3AvyvXHnFXauN1KJaOXYSovHd2cbA6EkVEAj5lCoWJrdViKxPOJtXch
sBqygK6VuwyLpmXIsSQbcwEX2AJQsNuoV9fQO9D8GmLMF3fAQLGGmcBRjcyN0lE4kHcB/C3JEBAw
wTYnAioXjLjH8iDizZ/TmyK5RQDlp+mm1Te4y8xXFSYK9ngtObKco4sxn/aOTFXS4wIhD9YTVKJ3
+fztWDAerNKbJhOXZixEaJeRamPxOQ0FNJE8bBPaegawqrHaSdj9JdhnxFifxAngaimyy4RD9IvH
Qq9MCWYuEax38CDlOUoVHV8KpT6s9tZfmeD37n4yWaJbDkXmmrrNNQcs4lOogR/9AQ2afbc5YTKY
2QuzlyJDGd7/aFoRWqt7fyEVKkR43fVh6g8C/jOBUbLHC32e3ipaghN67KSDJoFnRxOpe9fZadXN
hlbunIKHVEsDnOVZPKSoqj0jb1ftDnGeIN7Utdv0qT9hh2QCm13zGj58FTr6UrFriwxXdoLfE7m3
XZ1Hc8LWHhzxdGoi0kaZgjl6Qm9RyVKx+EhPMETApT3KhO2ZyprZpM9zvu6qcjInrCJE7km4+CQc
24iOIEPZMaNefkhfEeAMZy93GayLgIecVfLtdkO6i1BS7YOQ7Odqu0y5JvC31tS7DMiw28HF3rA/
kB+tIdBjFk8ZpHKUtuQHciXstpKXzJ3AkrRXa74KkRuxb5JlEVoHcp6fnKJvf49Xse+S/W5eG4jg
kX/ynvpbPns7jpZL33dJuXjZcqfUeWzoxdhMvfBV8UXZtaCrdnLQK6nkQfSUWkIkB2COLkcjTxWo
pMiBCBrZtI5nEWw3HSNxCcII0Rb2LeMK6B6E0heVX4U0DHkfW1ag/52gTjTSecTX6hzHs4jQuYmX
XHG4fqzIFRcVVNNgcLGpRBAnxqYNvsiOEn6n0Sv+lk4soODYkDeYQhA/NqU2FOObNkQEgX1MBpyL
pkutytoQ9cGpHx58SlD4e4h7puXImjz/a4RqNG/D/9d9Zv5aDys2OpqZLml66Lrh5sz/gNa+cqz+
y811pZsuvaSUJaMbRmQq04bueMTN1iEgB2eoNcJvXhpiAPoSGplNP2wvu/EJzlMmf1jMxysN6vgB
jqjWCT0CN1zjqZ4KNjIu7GrHf27+iA3D2kVkOxjD2pEk8EFwkxKsl4wRRjDgXmoOGsyw1uB4Jw5H
zRt59fuCLBBZVrO82qir/1QTisrbSdmZF87pxAJj1NhXGxdfOMzQL4IGubQnszJobRtEEQjl+Kop
tBzeIceo5Nfdqb3mpK+sMjLS5AVjyaV0k7mQrSeXXdr6mLBH2N9EdT0dHlNTxge/6+QRHC5jkfxQ
/NhdLZa1ZTHqVQfDZmH50LmRtYSBzo4p2FTKyJuvMeMB11Y3csTJmMVJxlMkyeyL5KCmkwqVkvdh
4jBjXBcJSYO9rS2nNK4xbMm4jdwUnYy8s4qFiwpSL74tzpmUHqZkLLuTKh/QvFpAUs7bm4LzjZNi
IYhQ5tKusD3au+Ow2S7qTn8Oe+iNQW4LoLHfyvnc1q9WfuFO1hxRubL3unQ3RDAnsK1Mb2EJvTkJ
/VydYa1RzsVeaYJ9KMnHzsjH8K1nm2M7YS17odNr7UPz9b1vIwJHCpsOiBSw2vmIQGIaEAI6BdQG
F/Gu4IDSgCeyO65TKlnVGH0j95sz61ZOsR73SFQNMzEpC9H8Ld1DEQRaqe2aZ3OZg32VbyCELYR4
3nkJrE6NkCA0/77+4lZfVlIZy47CT0jHnMyzHQ++xFuzLE9BjoQ6kJ4M+WamzDkgfgz+sfloELi2
IakCeLPB1o5rS1Wz+bIkRahQxjGRMXWx58G97DNhxqaqxlxBYWxjbVq3tdKAXjMi7UqKlIacGduz
AxOOI120rmYEmY8Qtk8H6jPtGTuE9mRODz4SjqdDZSCNtsMyGyVqMM6oFjPb36WLu/YsO7EREcBU
mYEiuEGYJBxV0tA7gHdQ+iH3HxK94odPZl/ytQAEXJHuhQgticjcdaVlluIXw1AAxFReK+utc+lD
wGqtpSo/uuyajvdt80mCmJPLEAzLGi1MOVsGnxF16tMKaG9Qkc9G6j6PQybOuzqA3KOZYQC91hmG
wL4kHrFtSN/S7YyjBtpgHbLSMpYCAsnZ38RVQo8PaNOphABzEVXo5CqsqSInu9ijDfLNZykWDxC/
kbvdHk7pzv2icUYMEt24UsfUaIAhgUNaq3KXUpDYC094eybjh2n/HRJkMRqC0g/PP+vmYxnjnbDR
vmKolp7S+AJ0E58wJZcNS621HqdOIlJ8JPCh0HvNwgHrFO74QU3Jy5mpCbF/xbOaBFY5h8BBTL93
Mo6rmhvRirLhShRRV69Y66f890yu+wkR45Nwdv6Jay5KtlKeMlWbLzQz2Hx042fNJfIiU+b2fcYU
TvtVOU5olHJxksBFOzCyULEqA+YHzL7X58WdtOAOeQXdfyF5Awkf6uSkN6RCxLAHpvtf4SI+QImm
jxjyrn6xitIz9FA13Ozjd1wfmV5nPaZEOh4Vk00UZFUQwUOgzDlANH6jLVoPZ/HYEh58Ikg3arSe
h6q/KiEoM8dVtDnmmW/CZNVxOPeq6JeEqSCJNn/oXeNTehEzjIZZ5PSzQjHebTQXMjAf6DbkqAQD
AqInDTWmjbbd/7As03YzKkRWCnp9DNx8a2MYEBHidO5b3h0LSMwar1dgHeF7Kz1b5xPiIQGLwE7A
wa4Fr/77e9C8SbufbDNKBZBAkAMVxFdauWAt3a2oO/vs8OLvB25mSObrI91F3fxhsY71Gi7opnR3
Z3TINny2Ztu31ro2gm+BcL88p0SPC7WNE9BtbOXq3BeyXPP2tqGxEi8J303i2NETc8LV1pccESxu
M6BBDyLQqO6ePNNa5P5GGKqtf7cnbtfvflS7NIGrpJxxIKnQVjpqy/odci3foxEFaxb0IPeU5SEm
a6OJakZ6kznqOBvHWLJ0ciSDcyXicqnta4D9wvxgEDX4qfLeuk8fI70o974JZ/CmINKC/ovPNJ/L
8PEnT7RsXUVwBeT9QI45oYQs+tO3n/gu/01Qt1FZNqw1h4O8IczqKDwwj1768k0qKDmn1V3n0r83
57x+axIyfBpxH6EZaxnxE2mS9gkE50LjrbQtJ8RDGTs1dabobnsUvOFIE1230oPkeAPQHvaBLGf9
NikTLEkkqPRdCQl0RobA2HH+dLBumU8xY6OxPqfRSBxNSiBWtprQUzp/lU61OJ4BDJ2t/2YAUcNM
C8dnvf0aQytabLLysfTMy4VPN58VGpt0E3rnMDirFsFDXXVvaos0wMXyq9mNkWVDBL2aUiyysWW9
OsMMVVGh+1rhFIj7ZwzhSuElFNwLHL61J3xyVVvb7sFvD3DoJsGAjh8UoImRWfZOe+SVa0UQJllz
eB5AjYty3QxCjIr1Lm6JL5dnY72QFPZ4iupRBdZCTHwuEucedtjGRIQLUJmZ2W/+qZyjqXYUl5kC
+8S8hYD7160CURFyeG1E50Ubp+zDskBw+JOoR1Q6O+5PLGbwxTMrvRCw8lJx6R3VgDWWlXJYcs4q
vHhatF2TB5X/BpRHqHAvwhLc/baCRIAc3nSAJ0dfVMEZCUth+OPDN164YUhac2blkmxuQU268ok7
6FpuHfIpR9WtV5iQ9JpMvYjfb0y1vliLIukVeKS70XbO/hHxcuZqUkB6naWVJJPLOAXbVEvverQq
lyc0VlohCHjAirNGAHLsAgORoTpmTlUjT3eFcCy1HzDEssosAMwKNO038N9j1AV707cCQb38YEau
6lrYFNo+4d8oUY/wfty7EksA0n10E2XSHtcFI/Zu4pCHiyGs9ZKq1jcohwX4/uB7MsK76dj1jhDZ
OVBGmAKOEHV8QkcpkX4jZNyxVBcaYhj210+EievdS2k4FX2ejGRecY5Go52DXYnSenFAfjJFd7so
mYimoGVh2IpyGkZAl/YNpqiNxFl5KVN3DiEY2eVEohJlc0+CpN5UM2DahjXbiPkb5sdWtVCJfnYs
pnA17ez4FIuH4e2+DdRtYU3vJA9UfjtCWe0iHiqjvnaBzmuoJqmj+yhipJIk+bohv0g6191QJYJx
Lr5wknn6Wenv6z0v+BemGc/sszdVmgocXnDnMIBe0epOl40FhBA2X32ebjOTTbFIgK2nGA3sDHQT
3Hwp9i4hXkU0HLluhaMALHtzY1t4qW4biTz7A7BCssGaJGxxHwx7kt0b/GEiEqpWo1UC6TQLEawT
NuMKFHobEehey1fWOd98sgYOX7dfc5Fl/2gmqjdQSh66OBykabkb6Tn0eiHlRR4EynWoegN30lWq
hJ/rWaH/fjZ49IzXN/vtvjtOd3uSB2VzxvjU/3KWbFpX2blgpg8z9XOUxEUmV4ACS40YOnaKOHDi
0f7/S9zg4m8345Gn+8GP03bWI91redKWdoiiW0A7lysFPd8XmZLLI0948Vyb7H7ZiLJ5QkxJLR8v
7GQJiXb3PdyJPWSf8r/88+3tbTAqxm8CjsSrl2Xx23EfK8dSNrt5grXURsvJSUWDYcI8eFOIJwaK
zQcD9eZbGRZw0+AXwJcQKjeHwlflZ+YNm/B5sr8r+LLOmRD0n/bMxKNdzXc0BFWJF7CQFPk8G5xv
Crk94dpVKkACi2O+nnzQY8m2cYsfCPu3k1zRcqmU/pAdn7IXZuA+VpXrUOeMifJEmFUUs8XWy/so
lJeMIXR/aq5pLKMR9qs14Wr7jScJ4QAAWLQqcJ00VVTzUjba5OvE95YXkr+iW2w0M14YV9sm9Ov2
CRfEOWx5vupvriGj3680RpxIvIVmvjRVxOBy4Kz42b0rIwsZHtVEH2xwEPUnp2YGE55VsNyhO38Y
G9DohkBcbPuttJrS+22SJdGmrQucxizcTapRYmxb3mliWwrxJDPZsU7vsDC71WvC2iu+gSPnvNPq
9QQB+gls1FB0RONwXiDgb1J8Ld9/vcbvHFVlQmBWlTK1vbks51YCOeNT4Jmo8AzcSBjWfWN15KAO
ADJ+di1z9ko0jDgocBmN4rnJvfZGAqj3rCb5TLCzc/FcDEXYd4faXVfYVI1a5BugaETd+1c0hsJ0
mCDBalSBH7ORAjKydDXfMKHy8dBLObIuXQK5Ydq5BIE4IHap8Lh8yF0w0b/R/9d4BwbKggY+JKZz
0MANh+ZYQrf1j8Li0ztHWAVKfkX9fNTmyMri3Nm92EqtXxFUB5ZQxGI1FODog1PP8afE1mCmGYfz
sws24OVdvi1S6yH1k8PqRuaqaNpJAk4qoS1fMv556TlLqobibDBQ6opn/3LovYFxcFjryxCFAzTz
BOyhzFwuKu1FUF30qf8+igBysFrLnjkGKs5KKx57uAqXz+QJUAnFm8/IUUk/C9EalmprzdZjNbbZ
/R1tWzK/udseGjyvnUC/LMUWNPsO4PEIRi4gfraE3DvSfSCW9zPltXp1vK01SA2TmKIcsHc9fTo5
AqciGo7MQS8z+KkWYj4QqdOe9Xk+djqoKv7EXEAINRhzsHjLaBabEx5+rWlkLkS4Bv2bv2OYVBAW
KzfNleOZBq+GZVFeR1e1mwZ0DS9uMdWPQ9kDG9kpqlv48/tF1jFJ0gVOtbDH5O74aWM70tszXKQD
k3HxlP+4KdoM7afNRwJHF2qVXYQ07Fke2ADxD4NqkXr0U7jN01dPddySrUEgSfe4X5BXBuS+7K4f
0eqOj8gAfzMyndJvSs0ZNPAfatfLPdxPaU7w0bFObhdmpXL8pN/on42CS00k0D4SCIEos4Q9ZPDc
nAjUqVbVfeybn/8Blo+DAh4EomyQdeNKdEteRCbracfxEYrGH3gBfTfa3FVcjVkPyC/nWauIoufv
du8bz2a66Fl5CbtZbxmeh/jU52G7owPEsRRkQp4WNXUgYd6Q6M32PQ+B6weOotA/8hwVdneHSto1
aG3kA4VPDK/XQkRHiIUYl++VWUTDlp82kBjAPJum7M6P7IcMYCNgN9fEfDyaw3UGPkyAeEr3r4G1
S00I2VqPNIAM2Cs51p/r9elBDXszWFtgtJiLtUW3LxlxCq60tdo1Jz1DlqPqxbLz3tvkejRsEudV
Aw/+JpBsDzMKcNbJqGUEBBPD/+j/uygoypbSi5DC1Zcb+qQwsHs09R/nh0/WzIGxeZphF2MceaJ8
Vcz9MVuFvR0SwX9AvY0woVfxbaDafmyk0r1i8mNLkocphgALwCpX+XyOM4HC8ZdnHQ74aWNwOijN
kx8usensn2ib70LKVkvMeiMy/Z9YxgOex2L5wO0X2PamHqetsweunrSrLfCwV7fOuDlexHstP7QK
b0EChb+ed6KzalUYYSb5CucbsNIsZODczx/2pQw5QnguJv2iAOkMp0BNfd7tfJmMSjr/woxVuzfI
sxnYO1AgSITJ03gTzrTAavshIWY5uD0KOXQCjj80vRGImkLE+LcexMDkJ926Jdzm9rHyStfQ3g8N
JR4i3bjFtNQul4rXFZeTQbHmx172lFIfyL6YlPyiAK+uO6UpzLyNltHm/u1TDVvvIiRAmo4OyXj9
Lj58BkpGi7lL+chYfd+cTtONkEFvcIfvJvKzCHcchT+R3Qo0mWTNttZfxKBaYT70Ap0iOyHkBj8m
/Evs+yj3exHj3uu00D9F+UqLD0/vy9OHI4YuyEmsBnOYqA3Dx4C3iHRcwd3a1jmTmVY9HgJnuSlP
0WkaBfplYOwWyxLV+UKQa5vBasaaS8+Z7vwOjFdR+e8AH4o5szEPWdeIOG36qlYqFXUlnqQA/5lq
eZfAtTolq8+OU4hSbctYHvpORj69YKFApUB6/Hsn0rlCEbXoFncpcK9VIr6UKN8btyx8vwkT/WOE
OqNDSmM4+bci3m72KMv8GyIkEmXu3rfjsn+GeptI7lwMuwfmx4DNVWtzwCDsHEiN51heI2GVX3TR
p/kUUsflRj9qJlRlDymooj2puo/4pUyTVoDGar6nONWrGPLU4cxiHJp/Jh/CKJVyR0/MO+bZx2Bx
0UM99AxkpULWGoKqT8F2ltZxgpQvRmjLIy9kxNiks/+jEyYI0fkytouC9scEMmBBuQwPEHHmMcoz
pf3ft6PJxpn9RR32SzMmW7WvSyWmX5F1DjBVFIkmFRN77ggEIAq+BEf5CQqFLH9IttMvShDpwIcG
2g+S+UlmWFXMEdnrSZM5lRcc+ImlAgqoTTX/AooXIdz1OD4MEfkfO0ijVE4+1P9gMrcUpMArcTky
qZiEZ8+v0AecJm2OKocbw88vhL1xhxs848iadutjpwQTaTxBARPlvPZ0KsjVSOdhKnYUlXHxSqVI
ZdbEBkgi0NnTMJ3eQtOAcdncgjkO+HmWRBChrQ7wzyeMSyZGxmikmATV6DpjpL1PhcwGZSNG8Z+A
j6mEYIRomM0/FSi/XLM02V640+5iM7wmOjd0yCtYqd0DFu0H7kO0aL73Rb8N19kFFwXrEAYZaYhT
Rqseh+/Pn6SHFeF/tnprunrKgzhpDjU5fD6USmOB9vRijdUrU9I+wJvqDzFmR4VE7pSKyPQ5wkfg
6YZCER3WZu7J2LBAffjdr2oxVxegj868998D6DS9iEDzdsRACEw3OALdyLLMnMwfx+dszTQRxcb8
fW8XlcM94NK1b9NsexLrpN1ICDUZCWiDdufEasAefAR82QJRfUrEDK185di859nMBmhMTNZv0ItJ
C1QgGNbl9iO5bM8eA2RX3scZXlDf5t2zCsGgJ4mf6CSSdtlt+Ph7PJGUL6tvAqvbMBqMHLivESji
pZvImHRCAZqY9+eRa0/1vUqJf4BxGsWANnMA2yWT5lvp2iJ2fY79f5kMoNVf2tTp4F1K76fxY2/4
YAVyEAJYEDQsVGT87WW/V1+vZZv9WbGi6pyU402tsuQbaWyy35ieZDCMeAjp527y37t291kLwlaA
myoEx2AcqS1Jj6IGYUeXr7vKBE3VzBWtwUDzPTtZ6K/v2VeOQ8IfThrI3lDLetfrseldiTGj/4JB
8DFfH49SdyKHSqMFSats/cuhlCK3aKDpR5xYCJT9eNHQwKy4LlECZW5KumBjgNFuoXj9B/aW0NRj
DOXw+bcvSfwcT7CqKdBMbt5xpCIKCZfc3Ppj6YnPglT2VsS4/5HjPt113Y3Qcyw7N+G1ILJGI9TL
58vZB9fJJMz8Ifv87MIqeWBfT85h4UmeKxfgP5UN1eWv27kq5J5ZazdmxOUUaSY3dvsHK60ZgOEc
cJFEgd4w/a0XarDEsCWAw91wPXIjrOh8qEuXLj6vXH7R7OUXXruRcEAv7ugs2P8FV6SvuG0uyfDm
QPLAiQmyrYNHBxmEdB/hba+MVTs8AxYWTSMHD4oPATAcVUXCyavonEMZijTtc0b5bxEHekBh2ocF
3zOMXreIV9CchYTngfzxiZiNsQrT8O5tqax7mVBKnP+8t4SF/itVejTp++YJ4mcz+JNUuwfuG5HY
D/l+W0rfkZuziwbg3h2giZIzo+aIH2wHWsKNyk8NkzKON1GVx/jR7hYBFFUQroeSkpdyyQxi+JI1
+0LLAXXmXI3Z7k0pNSU74Y9dUARk6ehHFpy1Y2ql/LPueZ6qJROIkd5h8tVGx4cl9igTzR52RkT2
iQzPfu+pKOEwgO5uSeGoX+y5++Cg726UU+24IEvJUxpgt3fvMbNe3lsCMdL+S86aHRd6okdrUmoB
fXBxsf3gYDX1Y7EA8dhaxtOFtXXcuKSj7l5f7g/WJKSuhOHgxt481o6S9PvLxzyjL7TnwP+Lxrfl
2i+8aoVjskVW6lSDiMwgrow8v2AcCdXcSCUgx5jqI3Owb+GZFsG/lfGIyH7TTg3jIRdYBahbi7MB
57EiPpMb0d0/cAwaSfxTBk6kdw4iglfPNcFqDS+SZ7Uu2KpBOkkyusUt0Ea/zL/QpCFkOLva5MJm
9E/iDW5XEVcej87J2I7+B75jXgPNwr6negvjeJHUPk6h0XgNEHEMsXzXKhWyU0Nx/I3f4zLu0J9A
CCu8mVWD+yioxEDiQC2HWUoSdp61VtrQSa3m8Cmnr3VvdhZOcHW27kIPCdsO1uYgkNunwcQaS7mn
EgRiNgh88VfIwYQPIvJjb6DAIAyPpUyZs3bjIolwMB//oPBsUHsALynBrAMeHdLVjZ83jV7Kq5aq
9dkvSsrUdPgpObn0pbHzMpp7d3Lmyp4o4fiS/mj6kumL4CdmMt97KbvqlY3t7qZZhbb0n0ToAg9K
DO82ssrsQJdkXUZWVuQavDEQmh/Dcnbz0ZKMitZslvjARMYEZtGvA5cxnRVxYa2RV3vhMyH4XjVg
X50hr77mzWgGuGvaZMHezbh0HUcKvZsVbtbbLEfB1zuzvLCvRY8f0RXpphOJ6YOM/VZtnowFWzKl
HCPFVTcn1VWVI5dvHxHkSPT8rk2vz5owXvJjFSX2GR2mcPkQ55Nzw7+dsduDHzV3l1sSyT0i17U9
fWRHDWE088XX0FUpv/Xn73e/WL0PH8qFbIA1qKHWhxN/FQGj8Qkpo1W7vud0sPu0VMtuHLXfenws
s0o1o+Ybssem/BAZpuVrmqEmen0L+yvbelqvjuvxlju84ccPD1tHXKQRPOU7QuQpNByXcZaSUgnf
EjwF3/v54wejEXN1kjVzFZqLyDXvc0JrYpElYxwZaEMQ60nU1kmc+ZkBRU/PD4Pv8uJTW4m/WNVe
U8IEskjH7cKOtJ0qRr0A/SxzSM6KbDNoeSON1Y4CVaM+onYctJrzrQzYoXPX2hXBg99JoSSdOyjp
D2m3AECtuJ4oJC0j02cX4MunX+sNFM3bZiDpqntprQb6WRmxG7RCdJ1CqhEqcp/tqnaunPfyt7Dc
s6lJIjs8pYknrr7QrIsbHuZ6+fGjCU2B1rDQeNakbzRCCb0rDoiT1O+tlQqXFcld9+b1uHbEyIrI
lblEQuftlSuKiASdsIXWb0qxzhEMIkbo4zP+H24/sPtntukOhbd3xS8ekea+pvBe00mBeteZ3oYA
958wQINOhdTpHCjqG0pMCPOekXanp0KLq10HB6bFm/ZHHwd18W7cd07p6GGjqa907D4XDYTCFDpX
CYeqOk1P9QcX08BG2kNFLMGQXqQnRA8KD+YqnMHF/nwljGbuCyeEw0A0fkwPb6Ucs4lepbrjnvE1
rk8Z+DwoaEv/NyX3gAPvSsy5E3UiJoBwNGtbc7AOjfB4YJ/aGZLacbCWS9rl2NjeumB86KgyoE8d
f8O3fj0ZEKjRD6V1MSSNBEM3FKYHP3TuQcNjYqTFVFzfivCrIhAg4dSeqdPihWIjMN+K6V2d/Uc0
5KQGA27NucxL+vtjL5OSunrTnbcFYRIVdoSFePZ/eyBr3j0PmgI5ukqiMe0rRPkCJPlPRewc8961
xGzPCcLgOTG7bh3tM05yltPYNdt7xVlh/StYDU5S8Q2BBHaFJsfmIhY9duK+QlnkYSy+7amGbWrZ
tbiteSd+g7NAPNUUsWtml8ov48TuCXvkH80lSOfzFDJRttHski2WiPlzx5GWtyyA4w+2VVlUcJ2T
9Z872p9K64I8DJ8uhSHdcvpkm4020+B04Gf+zi+9z1o+12uhmX/TINONsmqq9qEjZp5fXOgut+Bp
tWVeME/FpwZdK0xcr9F6twuutWxPWZGzB7nxChWMqnHJA4VNHhLdOg+Z6EGXxr7S0OS0gewKgTEV
HngOnVgMce8GbBUVs/22d5P9J2mxFBqe8b6h+v3fjVZjRvMHc5gFFOFfamBPRyzwApXXNgSz4LS7
N65zE6ZJhTKAJMyX40xCKQPFRevAPKgZFkASz5LeK7dJZZedZzI31wttfZBfCY+LIXYtPlQGcBcp
J2qdySGfXNXz5Wt/0scHgxw3rXCexBJjAL2ejNf/pHAFASARJitfOAt/8ohEn4TgzAWsK5TsHqF8
gha+17PRg/ict3sOqVOPH9Ue9nqvF5LxBMAh357gakM8IWg+RbIlG+eRn3XsHQ7PYc8phKxpvGtu
SjGgYCodU+ULkai+Il2fjxN0hdH63ElwIsIM8cpuJXNELaGv3ZoPM+nHw9XPcuh8Bv3Rt2XZO1uY
gp93DMrZ1iMQaGel6ZV0QunuEXXcAKN5MuwO2SpEvqXgF42gwbrrq9gaLZoThD/Ie37otnHxsxfY
CZuaoys1hkaEvcW6XLSnbt4YoHEG4kpf+vQNnAZ4WI8J4pz3LKH+rBgJQ9pivihKIBpdr9TIA3Q5
zsgNxHLXw7VX7LT+5im9xWMyRV5cGXeRM3JIjnuJXrR7hUyWi9NK3hnpYBBSH8Gq0t/XJ9F+kriw
DwQ7EvqxnOi2Yed5mz4Vt4Mui4MOKCR883GczJ9nT5qiVA2TUt2n/7GO6XMydHgZl1vpNu3NKIjd
xeGpqpiCPLbYlecpBQQqtIlXk/lpVR9WVClydj36JJj+YhjRPIkxepOG/6hZSRYh7MK6GWz0Yll3
NbZ5XrmNkX+3pH8gphn8eINIrswUm/VTc3z7NJdVXlBWpYrPOfUzcd4mjqK7o0knMP5QswFoe7v+
x0f9l07OIxoMbQ0dWlY2mzTam6sYR0mWYhlU9SLQooVLWP8ueGL2Yl0odU+li7uT0YFJLUFpmFrx
Y/YFFywgza0A5Gt6tu61WT1Tb0d+HEM+xayRkm24T/OfBltnYozrbRuYdrUjP29qvQ3w92ed1Sjp
74f3Lqu/wS4Rlz39iAWc49qtwVwPrznIrIHpPVY7K7CcETW4y84X1li5i2NezqIaa8n6fholhBwq
9Y/ir/HJIF/ekXtckT7A4DOJ8IhgyQBkBuLUpBE1CqdEr5Mzdc1hvifg6pP8mvDU1VMdyrybB9ot
pPLKduDV4g//JgQcd6CHdms/AH4zFGtJv0fwUV2IGhXefZ1KfGP7uYXWZI1+tRmwASDZnbcTlKQS
w8w5QBvWtce8I6pQKUn5umP5tfVGd4X/W4PczvMAaaYmRcOXdZ38YMZ7LQhJ/ZSDmH90/fZjKOAp
fq6dpt/IilPn+o+9De1oUDPxLFxZBHHdp5IUcd331OAbThUMxw8fMbcaeTrddgDikwgnaGatQII3
48D+KO/j8XN+ttvnYZjr4iehmBzBMMHYnZwcC+e6ldzqSNDDqnf50rmUKKZN3rBCVwSntY8Xwqet
12Qs0ck+4xroqdM2x/WU+HpS1jQl9uJ2gYl7kM4axCbEsLdSe3n10vtKngy19BqqrkQWt7buJjMy
9UByC2YVJnl2PZ50OQgsNdHC6GnwPV9USwMGQEDri08ES+0HpvgUvYiQA75rZtV/A11zpguKimtA
WQ5vh9a//8xH+vJzW4gvi+AkG/qgX90lIetMyXleuy/O+J4a/YJZtLJAFNdsXDr4VKQQI75Jyah4
vWfUEYGQIHw66lPGiRQ/bl9kJN84xgQo42ppcOnUeKZs7LbY5uwnvBWZF6xJCNAcxcVRE1x3Zqn6
dkV/qYlqem014Mi+T/lzs9aOQSF0A1lIV8y4AANL28dsx0doYViK5Hxb586uR58QZFqu/rMmF0jr
BuY+b0ppFwt2T3AZp+vltfjj6lcKKOwD4oKxdQ6d5tM4XRNPjf391NDLppHaazyCHHMpK/nBYWmc
CjZvsChekSGpIXrn/qPkgcrmWV5unMrXUOeL9yfgQ+48tR7SxKjEFN2aJzH6TnHJXzisgpAs4nzE
AYffd0V4TX8kEb3l1m+CUr+FnUdtyZvfzZY8yoYUGO+U89BClYfKlbaxVikG5aDPMeM27QKeMxgA
L3rbg4ZTgigNeuQ9wPpKsoBKpbYlve1UfMBBnsYMj048t9q+wtTPMdCmbPoLj37yHe+MY0RIEq8e
9A8/5/UmcK3pgA1TvUpoMmgjpwovXWLkTFx8Rj/vXbjelKkSGk/UzmClfpX1cytZlHCCZCljeJJr
BP299T/ijNLNoW7oDF2MxZk7xCQ2+SEv3asXDzXZXWSzkcyszOveNNsXqAa6cHOAmfyj7DqAVjJ7
7O1ezq0gi61yNgwYhoHHeyt++fYLBgZJYL2pRDX/QU7xgvxDCvmahsM3Mh60aPNoZTrUKdkcvV4r
A1AEg1DeQjYPiNLp12TbJ4XJSnVNf0dAY0Fg+0g8LhA5BszNTOvb8rMlfJ0rwhEq6eP8CxNG9VM6
5jNze3RlkaGzjqRc9uoVZW3pdV7tH6lpZIiIkYkLeID/9U92SZKGDiktoN7QUfnNfkagi1NvLAwm
PB+w8gGhNHcmXCCGhewGFvWCT/xapL/4FVOMjns32F4tx72Wo9xumbjSohVvSQj+vrH+KYQNpIug
WjpGOTSfylU9WBY8jC+kSbShAfyYum2zu/GYvEdXdeQOBEOumvxtrgDzBCIT5S6I0yzH/zeleYsX
rESO2WwY6NOaDslPUp9VvRTqjVW7jXKBtpTEaxmvDknv5Kqroa2NsFKCaQI4t0of9erMclrUegsT
y26zkV7OOfAtadshx7ZqfwNzHexvRcREEXdG03xffz8GPdl9TLSHnwRWkNjgxRkQ57rocTBj0lN3
4wGZ65BCWux61WM7j+W9DVYlepYfC+tbBVjxKyNfRIvcwB6T0KplYYptITLNctTWkGQJhTp4Vfm+
XoROx/T+2cAVthQlTC7nPkPb+Nfagbiq8k4bdZ4pZZt14auK7NrJFf6wOlg+8SQdKzsWLhLQv9Yx
QUEHlALF/+9AgonSQfiBuntG+tnnmI95gPymDMXd4gKoOZC1oA/9IjBtZ/hHns0Pncj4elxR7IBg
rN9WtuGnrmOZFel7b1Q71omQDn5nRUX6946oAYqlus2ZbYihxzAV1WQ9KgzmpbjP3a2lEnx+2pzZ
OeDZFFXGUSZZLuwCLFtWkBoZIvS4FanRR1ccAzkbh3+tlwcd1HKNUvTb/Pg7lfKoRMulgkq11iDH
ILwFjGlf9chP/Dy1rmN4om+/XbGBw2fWrzTLD+HD22hyFL/mwioCcntS5DZAB/ndsZX4nug0hGR8
fXBFG+YSyUOa3axlZPVIMkYl83RbkNBGKWG4EoW1VwlM2ytIq4Uh0sDmXuJ1frGfCf+LYI+Bll3R
8iQ3vJ40ZM8erL83xidLpX0m2YfM44go+V27reZ9x/VGKsBuMC7Uj+myR4FCj9+NW5wZNaRU37tj
LH+mIEABTjB64BkAR7OY2q2HTAWvVfB2CnWIBKjI665QunEL8Y/18bV6k9TmTioKcMa/18bWtBOJ
YxOxIqkYwr4umz918BV1qPkp3kC0+RO1WVyNQ7YV5EFMFFOOthWGKA3+O+3yd4suK8CLLy+5ZdsK
LlGROfRzLWk5EYetcel5/PyR2JuetMGLHK8WIsc5/fBxL0xFPTWm8xFE1011SNkCaHbNV6KyfDzQ
4vKy3Aa58+nEPKrclBME2aRM41WBwLN+wcGhbjyIdYa5A7wJF8GiOFuCC1Vk4iY57tWzpVP4ngCI
L+/mpJn9jh2/SsE9ESxFbFFL2wGdaAw3rD7QHP2o6m6jXnjxxhDUnnWmm9zCbzPr+zinppFH4G3t
EvSPSYu4zp2PlTJgQhHqI7evYIQHUabOiLrSezR0b7Q8cIOCvWr4X9naEglNVqskUuJTyVpOHdHK
E9sCYDoPk9yU2LnwyvD4IOyE+A3BRSTPdOPsElGwLRkKotrH6ebRM+8dgmedSDpCMi8ONrHVyKdI
EgTI+qY0mzNISCwzihB82LIe77uwmgkoOA4Uw0u7qGfhy6Oyk0+90FzLW9Ec8/yyxzaSpYfjREVB
aNqpsqOF3cD17HTtK3ygrCIEwgYDxqboUD3RvUu/rd+TrdNdxoR8NnW+j9iYOGDvBSWK+bxBgC6m
A+pNqbiKvXsL0Gy3nhxl7zAdZSCzPFM2nuHUbwl2vuugxc7pMhJp8V6EPRv12hY+stkiXi0Tas5g
fyRrfe/DZQmSeyKPUNw6dBYJaI5ZwwPA/py58gHw8LzS5oRLXhlHLSWQBRf3wuZJUIfw7jpgKuoh
NfJuuZYxQOfn8seRq0rmRC8BYj+Z1A17GASclWo6LaffnQk92JpTDwbpXuriSkMKb3TRT5IFfpJu
A5c5FNbhgyjfglC03dIk6ZFtlOmLRgDFhlDB+5jPLTwwIY1lfZd5+VqtRIf+it9tJ/7mmRBKpU33
hQQndso0AdI5jpqN4aQL05SFCV5IjCOGhILb3G8KI2bz5UDFf6nMMOqTok+ubQKk/mBPVACYXnV2
KieBVa2cvgiFnV7/doER+Ddhu8rxcsq7o6qIyAiK/kmdJv5lnhvYeRJ4SHU1facYknUpHCXG34iF
S6PGG9lakCG0qLVMKs1tL8WpdVXpZ8IZxO+f/poPpMa50zhHi1E01lnEPmw3L3+97ZL9nJjphRGp
blDYaIdQmnvM9Mz1HLEgF5mXA4fhJB8+lPxUwxUdjMmvo94Z0CbsMDwxBqzk2DX38HhXP1+gSgqI
z4BtKWugVMisf16Mb6pEQ0XzhpOQBfnKeg/gssMnH8Yh+h3YqxtPr6mDvlZMslK7bzB38//Oo9Id
15hIc6wrdRAHQsRAqCM7woWMGSKXndwv5yfUNxfeNNOeJq2CBwDgEcjL/MOzpifqIMgFJJ24lU/x
dtmuqxGaVeX5byT+YlY4YPes7zMPLkPFIlE8WZ//pGojwwwqBfqc1GxuXrPKk07M0v4REeq69DsC
nIRN+Gyj/U3U1OZg+WSbOVkWldlDZJHtrY5SsuFwz+CqSnOxgAIbvR3JUsGzPaHrV5rclkGfQDKV
j7VhaVBtA/BvyBXHp+WLdYYGcPQ6fckxJhI4xTs6hHkyKhPV9wqd+iKx0yFsIG+jWu9kdT0N1w0F
tofymvZhs6mfwNx5it8pdCK9O3CLvDDNI+JgcD3Nf45hW/Zy1cyIPdepM1ZlqQ1exlh4QOWALWh6
BHye7fwvsgzQh90gqTYFW43jquVL6GseCZV2PTputUuAAdeqRQY02bc49ZRTmmYZkjpXWfRNfYA8
KsSDL6nhBIvOM7wGhSngLt24Bm6Hhe+MH32PyK+fM2F8wJtuzazIy2q3hQP3HWXHFFs5uV6OoaIC
i3TGIQ/XhV5Cwejowi1q1l9wTgPlk94KCGOKcoO0WhZMjUbklaXJ2f0cOdU78B3sNNudfZPrHSIg
fUKSaiKCHwbvDeWSsd9UuPeU4wuN3bB/8OTuk3CjswY56dY//OSxJK/PCqg7wieIp8ypb80CNdLv
AH25M/0DlV3gBoz6O+nEpmShkd3zwzdOgbxb4BI3/wxz1P7UcDQl6LRAFf8eqOCuFbtCTwOzYftt
aK6X3sfXbbBl3tzHu434FNmqW8xjabmZFCB6OxfvLYiiB1FplPXht8D503CgLrBHs9g3tJpUaMO9
LQi2+l3t1WyQ51zx0PK80neAWhN1pIITfI6XLjAC7nGsYQnuYh3JeKSNDWxp1xzlP1QIsTRX1ctN
+BqMEtn6svwdgacXL3attRrhUa8mRqGriVYM+8LGazYieKtpCVfrZgj9CNFzQOu2/HArjevrAsLj
OMrM+RO1gHVFc8bS1ARUuiMJUixSUPduupa2g4+90bETr/U+dTZ21WFIgSdcUpwr9avcgPFruef9
N6UOoA7EyyrVdIviWriWHb4jRWfhIgrLNmCr03WjtCE9ILjlQrbddE/iVrtX9SaNGwLT/YaMk8Rg
enL828GPfcCxCyjhCIdlIm4UThJlCCrG/vhXBRxcVcPW/TvffMX1ataKxTGK0IwHBHY0Lr/N0oKO
jK5OcIurigawRUqdiz1lS0t1hgtRuj1UZQxURi1H2YKhc6Bmc+QFl3USqb3KQacYS/a64I/WSLTW
qx7Tb/gFebcuN/CZurRJWk/NCs+Lg2JIHh4miNHMNeMsoLWElj+fImjiWK2FutTE1bdObwZkIBRD
HLzT6zc+jjFb/sgOBQQ/O0eJ2f0Z+GYMJx0Mmn5uUai5GQ6/U99ZU8pibSyzKuqURoFIChZLHVWa
fO+nz9Fk8f0lhMmv09tfnj+sGV2ibAG3RrPkojlGk2Ua6WyEMyD3XC94oOEUCjSyHRe5zwxEGIxw
saRyZt5lq+KbTsu5+8xzZlujGA/TW0auDOFTFVAwJyF0ZWi6IpKJ7TH+/8g3VEGfXxGNIQw8hjFM
9JibCj7jNJ3Pcx80uW1U1/0DildmWxHVAnfjFOWOGe8uKahm7bjp6p2YGC2C7jV6KIzI9TJWOz7z
4zASRGxdgBXIfBKWD9gWy3woA0w8HKbWqkaywW7tkZwYbY9YZ1GGVMcHWFDtmT/U4P9LXSB9d0tK
OspM+EZDvPiB0powircgObs7RXikF5aKZi7XN8eVTsYWVMwG5HSaffyfJ3n6TwOB+8RDygu41kTf
ds4bwPpITDCW8oKk4xmD5TqrOTSgXDj2b/qgUVYPCZ2+6dM9QkdfvioIRK0YlgGU1dRFnxsHhdwF
FDiLxyW9yxQHb2lpyZ3GLvVAISh9ZcnYN2MBF3NLCrndYVCjA1y8maUTAcow/cfXezB8XBIwFL+5
zZ9KcvfiFnpt/RPLm/nNFjH1gCiOBCBWY3NqY63ob28v7C9IKfBZh0HQ5TxUEPy5lUHC1GG9A6RM
rTI/FfIyxAsaGvNq62AhNtK6aPCfq+SkHP6/kQ3Ep+66nRMyrmzedLZtRoHAG7UJ2iUu2j1Ab9HR
JfrQPr7NmTQzGk/EBLLdlGy0lTIyzvU54pGemELuTXSb0qofDItUGTv7zrY8ofUHVejwJ4g1JGvJ
CvU4UZi/Xkbj+PJXw6rnJgQWspExxRhAsPTvW1pUGW5SFFgHiSXcwGF4IZNBUKS7NNLaszsG9dJm
0qNBCLEg6BqDsAWdriaLn+nJSaP9LffYn8MygSNKO1C0AH6kWMu9nP4XdLI9yyESLPUbgFKyqFik
FsRqI3x0ZSl/SS0O70SY+8um2JJvVcBKKCByd5C7EKYR7iadKNyhYHQaLb+9QQTt2tot3f7zOwCf
8lJztmjy9cEm53rqjxc3Mu1GQEFgkw7ZOtIoE+tgYS5zfMNaVM0407Tf/NnIPDfImPfSvgh5rcUG
7o3hNJR0e7odC1XRJp142ez3lKe3rWBVg1a71WFqzhyYIVYj2f387BaA7ONLshAp9ifYSe2YjWwh
padg6lRZXXmg/q/hwYZoDqpzOnfhrU7O0AQNcUn0vVyWyviMqUOM67cDifyiT9HiLRGQK/OukGAv
vjAoYEEAX2t7M9JW89O5Wbe48Cga6t5IN5+1x0zrwqpshjbUOde/sGNoiKSqtQpOhptHbqaq2t7B
XUNlVVrohatvEOsvsIQkzbbEsOMIPJRYgTs4XnywUboCdw6GtIQhH3N1jWQ/rEqgQqfnn68nBuim
mWiJekxjXQnXgOBpyvgim1D7aoQUdskGjYnDAB+7cqrt2gAxfQOcaOIYGLJqoH3sNJWp12yHg8RN
UZMTbNE7E714bO8ec0pGzoJ1sLYPzhoJ9+xelbClsd4xsp+V+e2FX0qsHJVcHFU2BDW4JrHkc1o+
hmtIf2t7edUlhhOLM5XzTIGgjGoT6LDpgOm+LZsOlfV1lISjgiqHc/pnOXv2JhitCI72w8OZH0y/
gG2EHQX717bQUIKZtqIF2UnaZRV4lAGmXtvhlq+oQ77IFAgvQCTmY90Nl7aYs2Ki89VhS9snqxxR
RwZR0tN8cFEWM9akEbSiwJ9lx/9T2yK/2seSacyWGjlGWfmI2pjIQXddWM4FfXfGt6XUiDm/MZRI
qhsSNZjEKkS+K9NlE2NWNxOj3xMsbrtJNVhbaiEFb7FIR710A1nQQLn5DUVAxshkmxlVMntgF0JQ
2RHQeOaYV7XVnU+AOPxiDisGp4Y80IKaGKREB+r5rBC4gYpWgRne5MppEFSYwEKsLCaR/ojnPqja
dLv9d/RIDXZX4aRrV2zSOy8CwDXns5MoXByv8aZLLX+vthzbK70EAkAKnUI9ndaf6DKReuJz4gns
hFVB07hb06FrfClw16GrH8GXWe8EAYDzTXtYiER13IftYE5me8wgFoa+9idPeyU7vDlpU0PLCp2X
EiM9/z/xChuE2ml0JOLDj/WkBCtHaYcd9AHsg1Nc17D5nHRFXtSLuvCxnq7qQU6CWjIMGa2nlqJE
AcvjaI59iZCRKBsLJNy1SFVnwkMVRMgFF17rOuHF5uI1QPxSA37/rGCQFKhmasR+HUDZDTkEKr/J
nnmnaxMKubA6HpJVraF6it++MZ2zy8b3IvfqxXFDCrq2FPojf7gqezG7RafJZC/OKncsplLFJIeN
VND/y4MiymmX+APFdjtJpZuksxW6ZtT2EM0umFfxpU9oYFVnN3DvuYISlHhHn03lF5CwhVqXkYxp
+8HoWYAMqkZzXEW3Op9bF8z98liIamIt3MyDpPCdEjRX6sh2arKOv1SweZbyaDa8nATW/vVDseLz
dOahzDCt90YP2c29et/OlgiCERGhgHJ/GDRE6SnDouuCGsbI+1l6Y4TrGEVoTDcqxRXtNOIvfPkB
l1E5ET9QK3wqOfdsYNNis9IsnLBDvFM7R+Fy3+EvZF04w3MT8iKBBSnf4csf+zdW1mzyb/pocp8C
fSi+P7U27RhL/VxUIWV7LbbXW64o1CfDpyNOYJJfbMAiTQ5yhcxsADt/vgMUN7VkVWI2lwtyKGHO
zPD6zyCMrFILfJMb5/cdc8vImCEZaEJm/zPm3JkGkkmU45n8ww7ySJOFaEcD4ONPvIvT8QRqYy0q
BA0UJ2QRZf5m7crFrj+zkpevaAuLKMOXO07V7HLAnRP4MZynWYGH9Chs2Bet7xFC2xzgZj9mjkrR
5aHyGDuNy8soZDQvfLusQpGWOlbrixysktGEbx+t8Wjry62mCht+I10fHo5cYJAkq5rqxqi+BXar
WwjR1ztb65LzMwAs86Jn0hvCxC441IKMj+L88KSJDMldqyuMgfa40rKirHfmszpRXnFOsDiDRUZE
Vjy70mOqKcfrIIrRMSmCBZJ+fdSaJNCvr6cvHeicfbG85HMmQlslh50e9oHkm9gZpgT6TXh3jGr4
lWnAV7mv9m3rUAXTrYJaZhDgqoeJubxXK9+767XFwYOHzNupgengI0dAxFz+1Ez9QpZf2CSKLMCJ
eGbJQggc464fnVaC4kWIZts6Y59ucHd1S27oRPqDSgUnBLvaQ963wHX5V0CSIoW4acRVD1d6A0dT
5oixG4kPUZLUbHNaJoQ0kIx5WbpC4NAs7nla4aV2ijrCCgSkOHMnkeN134rkUQMvzrPNWet3JVq+
19WwOYdgzlNiQ/FJFZTuvpgttibiwWFiog2Z7JIvCVXE+sdRvBlEDQEKWc8pHlg8ElK5vn9EurJr
mPOotBBxZRaFS7VDfZ+VS4lOfBoNQSGvo8gWbLB5ytem4Is7CiWMZ+VvQu1ZnzTGz/8kTsCY65a1
N8682CDCdLNyey1ASmDchc9+YVapvIsnmmbOvpCrQH+lf3CaiYVPcdLMS3gOv/PRH8fdBWDjVKTr
Uh10+Lxl048mtsXpHiMmTmYkpTSIw8faeydWSbHZ1lKsC+tjWFpoNeU6wZ16MQ7EoFD2vtaebdQq
KAz/dEzU13I6pXigMxo9jSpaqi3vUoha+aiNVCB+Ff+YES6hPTE+94D+J4p9k6RIjRMJSmjoyB6X
4fC9rAD7LnAUkddg98AJgEpWFk3X5Kg30nI1OgNeO4bHnbFh650qE8mwgVa6Zp3oQha6MmxY1BQ5
EhtQIXmZL+LT/LTQ+fC+9K7BLAFcO7VZaHwHs6wVmbmKhGSnw+kjOmGXHsuqChZ6aNMKXlu+cAp+
JQ2ukKu6pTcW9oRowTXRYOeHdijppZN/yCaCMy4wjwPZrH5RQy9NHhUmfj/QHuzhfhbCT3tRkyxO
0EeofVz3nzdF8xS6utySQFtuZvRrlW771Xb9J8SlPMSRSiOUOBY2y/sf0b+qPh6pdriYf97pKD6A
M6tcCIP7+dhaeeg0p6LoxCGZrJTea2Jzxcb5edsTQKg+v/KkB/xaxBGn++EavnEFP6fEuLMhGogK
zsAj48/7EDEg8BcPClP51mGU85Tp/rtugRZ1M8fEwG0JqtzvMu6c048Hq5BgrPQUdavvGqz2qAad
2SQ+VqoTjlhFVZDEfgE0UDGkxhFGHNMvPnIAqf6NS6etSm/b73+2/9G/6paArsfwuoNjfm91+ei4
9hOOPqhHFW7hgQgEw/5JFldn3MPjnTlfztEbQNJiguT0OP45L79J3uhSmeiEaKAzifz2VigJgwHZ
mS/MSPBTddhnJsB40MZSYYQ/zUX1U0OSEFU+xhRZCxcXBp6diHVvLG5M8HOpi8empvqJmoOsT/F/
z4ie0yZ/UryEwrMoQhcY9PrFIhjiPBfJ4d4kPk56kJsmkAb6boiRuphZ/0J5xRKdcuav+G5ZblrG
KDlqzEUmxQDvs/pJ9x/pxwzYlE9YA2aPdbzGZJ85m+xl3+oAbYm1jMfCMpkEmhqHjk0lByWON6WF
rn9xueiMqlO4hnZXbvPntP7ezD91PifkKcT0+KHqhDcyCSytSQ2sJnT7VetVRcJgFcJd1DdsQipE
hhQA96b6mnouFwx+VYE9rPEkU1vmkKRScczgMGRSZH1L7yQ64BGF9+KtaJ1rf9fJWM1DTUDclcGi
QrJ7mTV/P++a/tciOeIGJYicLLbpGaGQbltV2Wr+VfADXGmmeTGkYvGLYNJM6FLgs6uVLhBy1GZr
0dxe+Skxm+vrvXDHX1ilXPfkFQ6+VHxFCZ8NMyMfHdK5vKjfIIrsPEMcj1fSGB1GR7KqIUt7rFKW
FEyG6NjEwJQ9VywLR+JAFn4rYyOosupBwhSdQQgIJLFFUnXckyGxklj5V2AKksOi388TKcF3KkyL
SoMgbwW9b3g8U6QbS0g4tDhCQ2IcPa/3gl3uRnPPWE4sEgXJZkFl1lPfkfkP/q6okFsOA49cmTKP
qEhk/BwI9Zy9mp9edrEvqLrKcxWJEJjjEClZGTePsNXeDtp/M+CKdqxd2dKSWr7jG1yzEkVnrFnH
hizMClzb2X19no+RKF2Gw0Jy7scVClOMZrzfaqgd/zFQdQYJKnKAAoEuTrKLZCTbd8XIJnnVfUFh
RvQDz7VkmFgnaIyGAtqO5BIMOwCLdX6bPDJ/MGLBx7udCQtv6juiBA3QTg7hpW3dDyLaIGBPx7s7
qTiXPSXX/4gh6///fBUJFMtni5wKAdy1BBA/LQlANHdugX2fimtHOyCOXZ78Rz509jSNANbcJGt/
C1PZXnlyu2vhDAwq7uP5NACwVRE6EMLpbTbBWUlf7vMiAR+6na62lwDmC+uLxiiSLoLs4lXnpsaT
6B19ckMZ+6ghFV0A+N5fy93oZ+nF23Yw4lugUxHXuBTj/XLXe+5Xv4m79kJLDLW/55GfDA0qKkTj
sleTnqIPaW8XFTddEkkgVZlMCwrLlGYtZi7wH77zxe3KwxTI9/73ISTBE+3F18Eja/r27zCOPY0Q
oUaqK9gsSTOddmPvcQ5NcjF5PF/zSxxbENLjA5b2LR1PgWQJ9jD9hYcHS0hLnOrcDVdu323K1rfl
YdD6///pzRJQMjmV6sJewd3GKcwChoy/q2PvV6YJhCA1YE1r5cg3DbuZIzGJe88eTmm/XW00s1EG
SMADdbsERN80ieyrM84yJ74KHaydQ/qGr3xPekjuujU/GvauKeMK7zAXkuWTNaJT+g+ysftItupv
z8KF+Qf1Q7Iij0df/YynU5f2hyDIbylp0nVJHiVQcpyiDnvC4APCHodPigdngwnMujgFdT1RUOt4
77ExxyIm87NlgH6cQqXkR/OBG1dOeLMQnI+W4jSerVzRp6akgUiLHQ6BZglEqMsSVvUtYDo+VXke
3ik0hlJbNcR5U6qLMRg/PXhpGQdhas4zJ0yjwl7m/xJdk/OimYrVFHcy1xC8iPfkT6Xy788Y2dm1
cBZBA1cNfdzQVvqrFIKuA4irz/eOf4wiBjewxcLXqdos3mGNOEUxGpgPOQ67g0cYT3QzvB1yonp9
YB4Vz82sD81+9pkDxK+Jo3kr64O+AT4fQ1XkPLSCPec1gAwmogWLrrCJUXDeA13DdvxLAk+Zt4VR
7HXzrllQyStUcQ/R6vRnUfUQKP4/BS5NLvv6xuBstOJjXEpFar9xfaYyxKQXsHnGp73boH5d2PQJ
Xdxrv4qfxHxOSpKpPSqQhLzqmBvQEawQbPucWyUEf4IQL395W8ZiKtWYD2RiGU2RWMan1ncLO23U
tLb13PgqK258iqP4KTJvg6mvzFdl4pumHnV7LNQY0v2L5Ucse+E10RYf3RTuuHJ8Ysyz8Kp/D8iZ
EdF2GZ4NAcYoDIknUhGDsOQC5mvzUGdI5tFRWCsj+HmAZdtjdinIBDEV0XJZkXMNdps5UbK4k65m
jnyiDenud9JR4s/1yuYpmhiu4fHRCoL9jJewEHsi6WXgls0UpTnpbxdjN+XR+hmJXtlkxOTeR+9m
QYNrjho15uQ8DDWQB5cfl71V/yLvu5JWtmPfuO/OEDQitzfZcmOfjClZcA7bJwBbsDqTEEJd9fQi
iEaqwZWAfe2/zzZWN3RRoIW5NWfYi9UV9+RD4+PpRozGjnM5deuh9aUMtLvP8vV5rY8OrySaa2MX
3T7aNCqnEJ/s+9DlxGZ7w3g9Bgv/FdwekKSjdcvlFf81GtsGGTb4h/reCpTUYVfHvigvk653spwx
SScE8D4EFLxLBFFnaz//hvFvxKkuv/Sycj7NYcepklTPbzYSZ8Npod1NDGOZ03NiN0a5VnbGnhc+
pyG7e7ZykTO0Uk73YMonnNzktxNn9dovWYVJqSBk+vUUwQSWTorQGPV0XdedepKbptVrglxK2tBX
zBTI51Lbipj5YEDxM25C61T2JaozzBWYgnooS2qJeDQYlftM/RzNOLvPgpxRoR0FWGRweEUcKP8C
XMp4UsrcgYGiZ+Vu+GR2n94kpgePGp/VZRiZa9J3I1BqWBsoOXOUPB0qnWbLe1K1sWR5wVdx/Cw0
o9ixSouGaOEA3PhIt9Qn90sYfz30DoY8vtYcp99tk/MDQndrPUJlOjG/yD3u85RHJ6mVOcTWJ3Sw
p7Mf8WETXujbYtY35mw2SBpmfzneT0O4fAEw+hoJsMzTTwhHFnlJBNANmF5brF3A4MKK3L+GopGX
v8IuDDWrJ0p0Ie4/Z4D/9ERFVR2DHr3wuwNx5u0CaXkrGQVMb/ElgyaCPmUlIwnD4uQfJRQI0kmK
aSQLzkIuU7GKAYA9WNo0/aLRiCnUOiBuuyadcpji40/YOQ4Jonu/sqkF7S+Zmod9AMPaD96s57Hb
hCvcocHZWTXML0AffzKvIPAKAoPp5GN3XMvo8LscyVEDJ0w11LZRqTo0hIQuLfWG+/X64eN2m8jg
Pxyn4djqaTvaid3eAD3K9JfMZtD9yrIjy8PvPh4ANCNMTm1pgO5Yz67kEY9CMDF9z+kZJZokEgF7
ZrCEML688HEwddqaZQR+OOrXLM1NlRiuhtyVf1t9czRrp4O6pC+Ak6msPis6Vh/PSM2zLz3fJ8wa
Zh351kQOE+eb2evhQLibaDiyzZrBbmAVKcv2qtlhLdcl1Dr96+ibg7b8t1TLDGKMKzjMSbQ/5UwK
PBHJpEy09n1lcU+krJFVq7IIR+hXACrTHmRCd49rPtUDSqzr24/tVQbZY1GHPkGFrMpcxfaOW7Id
ajzpXSx3vAXFSGf9nBsuVjPmoFYSlsASWuKnwE/0j2R8WjPyh+lBm4vO1bJPJtHufJIn6XLaio6z
Kinj+udUU3V9ejB+ebYxkzw//zPA1kbb0CuMOAIVcxdxA9rbLZO8vQl2rk1CMCAQ+bBGlcewF7/R
8Cf/eE9l8LC9qcMU02cftckpt7F1bAHJMEOsVIalB6/PFDbNog+mZ5pMAkSuAvgneRQDEFDlcmF4
0stsyXHNbYa+omRAtIJhnrv71Qor542+ajIEm4jy9izTFfowkIPr9iGPUTQTtLuCCVGVnxR1HMMm
OXUxL5JuCJZfyaJi8nNviiLzJe9KmEYl05d6j2L70TJt2WlP6TYSl9DuL9BKPmVkKUCJVWx6Mfsj
U7XHSoXbZbyZJh5sx5DpTqUinsIiCQS83earcdcCpKPIuYJtOA0EViPUw8v8CozX44ckD5jVj5eb
GdSyDVB5OucA2rVUbMN3dH9gVzfRiCoDBbStt2CjUhwSQhbvi147cURVA9tNld8wjfAK/q55l8Fs
p95Y5Nde3BOAryRQuWcwjFUCjLEWkIgsgWMmiamuamrw9TuzjOb2vcNNWtdMkM9MCY8x4ne9dkK2
LQrfFVS5pAvM9hkiBgXhv57acTN+py5XhCo/fhlcWg/aINfHXzQBVzJ4hwCk2YknCUtgnkeSIooB
Evoyye73uFTScob9XTgNExIJlJVdv2jp3aUdgvWwu4vNM0MrHZbl2Ci/hEkWOnDqjGxaAw3DycCs
zAFmLbtCo4pUVllSg8QSfi9YH8R9SfTDrdAkmv5N2W19NoRNJOI9cBR/nYrVIwoJZbpktHT8aLrr
iKnrEkCxiXYkCxp5Lm5LuZYFT5nMUx1wxav+SFHDX06W9fq8efDjuqpCaAZ9LLKeNjX7g7a7C1L/
ndul8KmpRdXI/hOwVa9+dnViCDCBtJOSAc2QKAv9NzHbcHrowIM+TjI/5Q1se54XyUte2Gd89Pc7
rNjbC67b4REgZV3wnoT4rGgj5BqkaKSs96EoZRZmUK5Rk0OPc5GPPgCR6+XfmdsjltmnxTtqOGUi
YPxbiUwJhAkJ0BBTJVsnrlsw3Z/9j+HA52e8hcFliYYiMrNjs/hjooIhUBS+BcjrL7QxWa/ku2wl
XwgGB6MahGLd6sDFAZ1LDDbgNHIgez2siAgx3K0nPHg10poAD+SuVGVSv8NgeQxIHdyTU5h+0b+0
HrG6hmdT3NOUBq25q7BstPO90tZ2iuJaMgrmXEzqXz2ia+ZZk0btz7q38KZ07RhAQ36KuJo7uYgI
A/4zJItUtT8ptSQGHec+lYZsHBYwSWgE0Q4Bx2gY2PNwZ5ysp6YVwJSQnm8SkrRtFSM5bRAz9ank
0+jrhqC3wDu2ncAIXNCMq7F3Ev98nCxt6XTc+F1097gmbtDPHnFah3FDvrdXZXmkns/yK+aIkjoa
+5IanTUhhD6d2pYH5SBaP39lODo4ONJ3FbSfkTWUUA6COLUI+OSm6Kkqs3J0GcQfbh2RGNaIdi7P
I5lhKZLb1AxHjiOZ8bExPb22/uS58oKMQilVRCGXZ/EoNGjVyyg1Am/XrImpheZ2x7YYvFdRgsl5
v8PAMKb0S7KPUEBQv4wLjEAOTpKwXjqJWhf955784c3w6kSuT492vBVSFzurVZuMFt74QTJ3rhez
vrHAObjHjmUNXN4oO9JCMCcUJAyNRWY+Cb4LOU2s4ZjjY3SedYrDjp96xo+poYmibuvMWohNGrHo
UzF0mEC2nXg+SKKbrsMK9cZTK9FztiSguMEVFhYn7J42m9CvnWcUZRZ73OuFhYam/AczDffy6Oxo
EsJU04aCcGfyx8FOauUN6vADP0GQIW/y8wdxo45AhFe4yWHhtf+jS3Q5OfZoTaZKr4ks2y8niKxZ
3MYP0s+dlccfHpZ/SQ9w/6ejY/mW/Mqvm6SbJ6LdF4siSHjnP47YLw3a2H9NNND7j8Wtm5Qv7gzR
dZIMVvXAB0fk81kUsBhfmhnyqlXN4MyjH/Tsj4t44zT6TTkPaNfNhghxaXgJiIc/dqhwO6/X55Z6
2vVZqOkKcc1xavMLYJ3Jog2Tgr+iYcO2jB8i10uXwT6eugdbuKC4N/orse5Z1RS535B4g6OR1wvL
Jt5MAGJ+cYzbTRm7pdyn8z8q/ayX+L4nonpRFvKs4S7+Y8Zrc3XQNMVFVvH6h/RoIx+9gnq3Pmoc
fl5dJEqjtAWFdQCsuQlZkyXyBomHAfPG9h0BW9C94jsD5yJVnAsogZMT9RwiJqX2zGa9pyV4BBe3
94ficfAQySkOpyjF/6rZPY0PO/U0NS+gjW28XDZLCgTJIM2Uwv/5V8LxjIP5fKetfl0cUI8kc4cE
1gtaDoFkxGG1Jv70Kqv68wfafTKtxCM5KcsY6Pk10u/dxl5dfMi8vO/JXRk+e4WYtHSLj/Uy3+vR
vSQf/e2pVEldWeQFv0ZMS8sMtNYhQMiTbdeNqYWPJg7DTW/OWaD9/R3Um0pUSrtRSCnlH7IHFt/M
e7fC1W4JJCL6bqCxCIL0AyCb3hQJ2yDwsgCW7DPoezOamgEq8dhb1ZOeokFOykDIQ9yzk38lvoL/
YZyNbehWM3j9yp/2pe2QbSHzZ1uPFtgABz2ZtDOrD3wF9VsefBfcKpDkwW2yMMKaG/7ZXobnc5jn
EUIgti3TdbU5c0ty6ihM4moFkw5exFp1SEB9Ul9RCGZJcj2/RA56PH7w75cLfT8KMHoWF1sAD2Ue
/NgzW6iFzUGpjkqEQ36hVq1Bu4iw/VXNCjb8Vk7VOZ4nLykXjVKDm0xgts9bllacmWwHKdp2UxQG
l5RB24J4RK1X+QUm58pcCn/8HYLxsQRG+5TOrLfueK+NxlEoN8Eh4ovJiFS+bSpInTbdDc4/87Es
+79X00VPGGmoQNWUPR8gBPzc//yhFfVvaTJusZlqZDFzOkKaVAEuJ+OsUazzGk7qM6Tkf9xErzKd
xmYaYxqdTSKJhPkMNI/ErILzKwJt1m5z2k57J6w6YvuKtYnIH6XXcoqEHXlPEaI0UxzVmJ0L6TmN
XGCtFCRqj4v1HOj0TCvjf5jjxq1aN7MM8+PLKdTC+E90UOodDhbsENbVR0YFYfXoVbWChpVxJZhN
/RSV+JgoyX3CeM8F+mrdCqBJBmlKx1qhtJ4KgQxfUE5+Gitwm09HkzRfSUKmJO9rz8QGaN20Y/bb
gnByBfwPqHZgmWZa1Gy2cJTUkyfw2chLs4UYwVUBjwqNwV9sEtt0AtJLdlQQTpamXh5B5TMxRf1l
3BR2a9pZqIB6QoP7q4huhy0XF336ZKHOy0MbYGsHeBf1OBYNYK9MOYUZgo0EvNBZ0u9TLZmEsja/
wDgNLtXwLUjPZi/g4ki655fLME2okD2OwRydWbVhC13CL3YDGK1S+pWOxauKMpCxM70mivW4U0/K
fgbFxpKM2231XvwOB5ZnhVp18e+4X/a8v056/FGGk7dR/Z+uy5ZT9Ao10WDm03gmex+GaaOWezIk
VO2QZlLeIaS2wsMVDFdD7qv7oh7nLDu3deasnhAYemk7nbmjMhHcpYfi8DW7MZw0vM5cjV+6vDBQ
8Y1IAe9dMxqjwooWyGTzdT9wWG4qsgOCcSYOcR0f7Do27erEdpyDy43k02A8nDAXAymM2qC4T8iw
mf3jCfdL6RucZ8Q4TtGpYFjzHq85a0iYTbmb9y/sV/9m09XGGvRNONhfwmia1gOLpp0RAHfrg0XS
ZFSvu0l/7eTw0jhHabkQcdJ8fT4Ga+oi6VchdGHW+WLtZkbA7th7Me3fFwh8XsfAtXuQSppFgt0b
x/ZnLUEzA/rAuhH77y3+LrwNC7FpIEKVUZECBMJM2jvOceNpEuykpiECfM4atgNQ2EjbPn7kFE8Y
5TqN2DWlj5PZ7gUbFPjS087Mvm7k/1tv5GE5TmOzvLa9IM5NBQ8fChjjqvZDERqjRMxrJes+UqUS
x7PtsZBf8TV3S6gm38yj96CRHlimpeppi8nQrAUIU1LEkosnwRl0YGvYuk6sDu3NMBlNAdvRgMe7
74+9dbIqOqvcT31Ou9shsn/VG2FSQWWctR7E/xdWYYqxCURv88oU2loZmJC6IkyYGTH75S+hAG3g
kx62XzYnXzhFNXTIi/E7oZucEx40lvCyCcJhXkow2/WnLKpvebrx6lXqYrUSAr/qhYGmrQ6nQ7DF
YG+t0A2YZJKA0ibCuGuxM+15Gx7oTf94naLd/+zwPm/G/Oxv/qWgrRarkNjzgDJBY0fuP/gVwgDZ
hZZ4cvHCtYSRuMGjZCfc1N0/CwSJsAgOIGtHD1qIPzw9cOXTw+L6lo61ziCZCMdlGJw9xRX0ofWa
2zu3Z3loTIHvBOfBFhG/vIknrsml+1sf/borVbdxxao79/cBTdRQTXeSOiykwxdE4nuf8Q47FPWz
oF54QE8ME0/QYNBIJLaFAhYNHyQpFF7rY5obD7xnvCZx8P07oRLDUBaMA/5i1+p8MSfMGxfCqvur
tNUgTMW3KcQ/ui8nWtO1ZKj/bZqvk7GzmCzFQK/7Kfgtj8uhR7hbXU61PoOXlFRQNn77y5ASfA6g
gw/GxCMdh2lRIBy4D6iITi9xsV36H7ZOQkFlN6oDYaZPKaOQ4VPn3nsVw8c8TU1jAGzKfkCyv3WB
/NUgy7a19Jyd677C8G6ACn6WGxWq8ZNPRVb0g9cUHW13Lj5p7wIWnfp5ME/lVsDMMl8qdHLNJfWj
hkKV3j/gVZTg9T6bAX1YYoF5IoWxsSNkt43gPqd9UPjLmIhpC0BQbFLX1B5KMQcPAbiqydEnkZ22
FAL9pa9ECF5VgSTQQdt9fdBEttGN6gw9BTteX0FYsrqLI6HL2pX6Ofc2qjaOrDLLFvT8KqkoxzcC
0YK7M+CD1JU8VhbEVWD5yKjlPj2/ryezPj4cjn9iUzrC4hJgxL4PgI0Izclle6kYmUHdhuJnoInJ
PoWF/2MbC+46WiglbA2w6U++79+bWnWvnNmPnwRWZtQVhFTWgulQ22O4pe+J/PYmBkKLZIcXhlDy
F9XeHRcU+KB9SjhJU7J/IRUbCgAhoWdtI1ZzyWwQx3ezP9UipLk05nR7YphEGByMTIrsW/JQowdP
F8mkv844FdLThc2Spn9A3J5Jz2sji0vFwDxivCqwguTRHxG5hqqbw+sitdeQzDsiCvcPmy3Fg0E9
y8VMUQqhvFK2NQIZSB+hzSSpb1cFBSOXxPP5QCEmqIseeOgZ4Steuz+mFxi9qScL8iJIyQyU/IGt
G9OwbkIVeZRYP6K+VUzvgopLV5EQCctTr+cmem5ZUbJzOs0+N8noXQyHVDWhXK0LVQxNhYLNLIb8
IZ0AvyGHp6LUjlbTQyYfahUt4MYxVfWoE39Y3ZYrfB7txfrek+1Q3nM5n+VTISgyajjtMY0P/8Zr
tSfwA4I/POfz1hLl0uB79VGOXv487BuyoFI6dNURd0BTEWTkn2LXDmDmzoz32rhIz+llrqUg4+v4
3fLrUiXBA/vI2N1Q3gdM0rUs92ATm6iDCEjYyjlRNAwaCrlrWlLzjGmrmxdGXxZu92kAxoNVC8mn
3I2fZ7zTHFUvEvrHSkY9Sfzs5TSnQ4lYjG0dfKGMAzgx1EjhKozk8fKQoT5kALkdePj0SO4WsYad
fKoMO5UgfPS/U0Iqcf0HFYM921iFYAxD6R7P1hoWhYM7otnWFlcXebszpE15UmSi/6fPOEutNOdD
fMOTMrqYQp+9wBDXSCbLfyTCr7mJ+JxpKxYIpuSYuCtE47q7RxiYCHLWU5kEOnh17QYvOmNfRVwR
N0Q/BgCwh4i3+V53XNkOJcm+kEroRmdP5b7TaVTv3+Nae18Lp7O7PRlQvUurV84KhOItCLeMpua8
tJskfw/K616MgsxS2NQ+Zm5HQQ3yFehH3MlS2GEmuS1zd2zOekHJbrWuZaM2P03pyAmNi6A4wCJP
bha2fIvM64wyqL2yCa14bBr2lfuH9PoPIDGPHRqmblszS/+ol2e1zfXboDxZ2dTtbzz+xcIWyEBX
gbM9eCqkmhkN4RVaGcS6FDtj8+lJjUwNoaRtXUj3beBKRQjooosKhXIa5CWWrMBqqTsy+orNuKLj
zb1yIyQWNCADaWExsMp8408qQ/cmJ/VGpVSLk/r0U7ossOEcffCl1her86yMtzJlA0UoB8x18icf
VbNMY/yCJffBoXhifRuCAr889KPhuvz8EGRR0HOaRhH/7CTW0VH0QXwsu/9JD8DH2fJ93Re2zvtu
NNsAY42cRxrHWMkvA7z62HggrVb+VR1JmkMjqX9T1PPrAUG7nyChoNNaiC5oari8WO3Cq9mZ8DzB
EbbyUHZ9vw1TvacIqvhpyc+xPwqXwSmOGRMiSr7XC4HDyaE313RE+7fEAKQXtdhpD3c/xyRP+7gT
amdefWYT/uULhH74PVc7UWh6l2th5iWJ+yIDp1Kui9LaIcas6ubsfB/m/Cagqf3CwFxaOzibp6Rr
UXUfL208bVxrrf5hKRi3NHgAiFqX6r8wxVZ0rK4xwMRaWUSPOml18IIMaDAn9BjlLg1/V6kDbser
T5pN1vfheR/RPAnqBe29SdoyXZ2g8KkrgEKvbU7oSzQ+CNYi9JvenGgEN+oCs//hQPxf/0ugq0SO
fsk3HtjBLJRiJOm2XEV3lWeO0aknle1qcfEikToAJE8ZFX9KytQohKqJe5PxYVfvQhgrJzMPHo2l
atd+jmLWJpELBKN1oEo3UcRCERS1PGSlq439sTYGBPHSbM2P6bYA6Q47PtBCJMdzcOOYZoc1xOAl
ccZoWMHgZsnTKAO4OHaznJwPmhvZiAwhSRGvXO3IDwkflb8TdZuDzfISr9TnEIa4F8agu2hbIlex
Y0ES8beVk8DxaqN4osvpDisLJMYBM28V7ypI8Qa29M5FbluV/wFx5vHTYUIBYGGW7oc5HGcMurUi
ZcmALa+l1G3Y7zCjeEX+BIeIV+UXoDHwu19xPabG/JAuGxbIynQgIfrwLhel+VglPt875Fujjjuu
iWMVJCpWnr2VLvnPGoX4wqRuVg/3DwDPbI6G4I034MkEACjMn2AV80sKRV8QxSPihExqWu9cDSe0
FxoSBqdiZWZ8OXvSjm4jAI5lxwxy/ESn+pMzSFIKkzxOs4p3NgiskFt+VFHAokhB9qVfGOwgDE9S
7J7QVkwZI2U6rz6R7g6Z7XQbtbxA+xAB+3I0ZwoQInDLZZqGNhSyhem6ohm/nm5g2sLo4GDQWMQl
IDg+j6Htfc9sVbObl8BvrxA7s/zcit2EVHl33OAQoGxcBl2tH17GyxNR7C1wm93C8qRSjQzxtcOv
jrmsUK+wvnZAjSRsNTbBo1crJA0+vvDAisrML5n4cFih/JG9IxEBMus4TlZp1zJOEKJYMOFak1Ej
hGo2vWKmnnu/ISGsbAqE8+/3By2rAsfoo9n1KAxpCgVOSF4qVVbl1b2VqHyjFwrP1s35fIGWH/v9
ha2JtlFnj0/hRZZU5QsEeugS0KWQSGOaAEgd0yFgpd+Fra6RICmKAoVqoNwuVqtvJa4NIH7OFJIg
7n8tr1tlJUi5vV/y6/oy9AOX7BtA7Vn92sWN6O2KRPBqMQfvA2kWdAxA9FawJYpVgkG9avYt3Q7a
j/dyCm7YHnXjkYiAC4ekxI+lIoINF2hzCOdRZsoXG3xHivFp/b3lGc29lt7+Z+t3q3ZsarIhAiK1
j3wMoECjx1SJQHcYaI7CT1DLurxObGJSKD+1No6F/23XV4UMZ3O7UAE/kVi9rDWn4wTWMjoP1ZkD
6MBUfYXZqLxQrleUk5yrvBHFk2wTa8b6nJcPdALFIBBPI5L4awWVpoVkkshaaURr3cTDSDVhP5/d
mHn8r7cWerSh/Oc8ZhXyfxFm5/c/b2B/PB5X7yfRNA30kVAdMJJA4nl1E+4Q7ky7J9ZromhlqiqF
aRjFeDTvFBum0vj8CovHccxgoY2eKj1020PpI9tmVdloXvKEyWsJxYH42PaTXWZw87Mr3tBrDIVT
Iq1U07k0cKag1lV7Rhb0C8AIPFn2EhbVf9xGhe8b1/W2lTUVVwL6MAA6furCuYwXqOnE0LxdZIDv
h110RD637pJTpMHyYSt8X01ES9xTU/VnqC4xElt3VPMvDzi+CO57sYdjJ/qshhn30VFMkGc5ze56
lmK4UL7sl6lT+ocvkfkno9SN4F/sN4JsWx3OfLDdY1qqg1tR5X2v68m08QtNqRbo5qi3uHxTK8OY
CskLnu37WtAMY+AvLIRrQrq4+U9M80fJK7Kf4eD87/3dFhTFFlB+7lJEMrcT3C9T4/5Z9Uv1eUCu
6Uw7XEzuwcdGFfbQY9JYsOZwfe7COsrFQBL1Ttw+oUxs0LUPDisczMiW0l+XPWy/v5jboZU6qJKc
W3rw0MGQF5RUrrM3tf45cxrBtmVCSJ+SB5OhFzqNsouFxDoQy+8f9DPbul3jffLcsiX8Kno1fDnS
ypC/3gk++MVZAthNtN59mF4Gxcm1q+6DnRLmcF4sUQARu6Tqkd2vMdlwwroqFNOz9pgwtIzutW/a
2WtVyU1wj1f2+dgGkgN0TNlpGY7WiphG421YYmOvhyqyic1adckAroHrbdvlc6uBgcBe6XrB05C3
+TmKtUBGolTByTv4xWnp3JbdSc/WqAYplBVANbZB0fjekprPQFKYN7W63f7EYqIKGJWRJb9J5Ajw
/zrPWALyF5H84qe3xQvF0o34s3BqtoPfZYRYS190ANBwsozRDMsWah0QpZjYPHi95L8N11uRtWUS
z0tkS8fbGMi+E2SDjQFGXwa6Qimgr54l0mm3oF3mBrLrz0rh2f7OI77/XqVEy4z7DKHei3uXVvYb
vD2Rt+Zgf0o8pBBPTnkD8grtHA9te7mLRASSJ6ETxQ6Of8LF/WaV1QYEz4MFgbUpwDQF7QZUBXaA
a+6GXxetiFpI694PNyDhzbV/8jOTm+EW7z+rdCsCVHv/0ZqcpjJTOdluLjvnpW8vtU95yP4VoJb9
+o2GPvs7pt0jikGpgmpr4j5HmkD+bdH3TApxDkNcFAt6P/nfBVKmJfFhYPyJRW9qhSwyyAOkXTgF
8SrxGoe1820KevHTiB0AM7TwXPDfUOyhVbXQKmswRqlBrgjMplE86o1xkigcyrppbXJFpDFV+Dw5
3noxSHeHFAt93wQRjOd9wpBVh9Ae2mhJP998JmohyYDBhQ/6jFb1n77XXWayJJSHECe5BUmZds88
nMn2rSy8rp5Kg9C9/StWgImuyDBnMwhI/BC/323YORp9L1WbboOv0Sjx+T5MkzOeHRl5Ty0aqu3s
Kq2NAl+ITcOQ5jhR31HJc9PfIBvHU5pZZPbljr4pEYxCYgOKRQaef5ZwDFf3FoE2Pvsa/H58zO+O
ImGpYl17KoprqGhAbGMjGniNCUPhXSnhBDrAkN+pFxiKG/pjy9quU63BYo6VwrrIugtkk8bulegw
ub3yfCb3BD8fW6kWq7r/AQm8vXuqOa4nn7R774e9G8zCSiqGZf/dwCIi+5LqYllPLuAyOudXpBd+
tQVmXnlWB25nXUU/7l3Q6cBwPiJGkzxEDlLn6M27aKpfrQMf4bAFdBdry+8vvKE8ALZtc2JN/DdM
qlvWNEPCvYNHuIvs3VrDfYYwuor7AfUThkRSKwqxExlFKMg6Gh19vMRndFwxuNotTjba9cSsYAdS
Lakxn28XM7Z2ft4Vzo0QkQHmQoLZ3VeMh2v+m4odyfsZ8LEDSl2r1l7iJQXG2By6TiOLN9rCY4id
JFah/DCW5WOwja4QV5xuFMTJOm96uo5QlLW9CDKeDpT80uYRpQvSKdoO+Y4KkSIhjAgEWJQvamfK
azp5urzRQeNeHb54ksNKxZI1JiNfGAo3XRg3Ava533EuAfi+XX/351f9e+6ttIAb7qlmjhSA47UH
OpGwMJpwQjcPtqQH08/At8mnNfpAvqfJvSGzA96i4cBZOyYoDbPIgzeGPajyUnnQlbiMuxgzKq8P
y2RXew4J3Li4a7fnP5a2bqY3hVaFj+RD6xXyyoUhJ8OAOrCLryNV3CcYbFJIzCTU8lHNRkSviqaV
EvUKgiRKozT+TcYHGCeRapaGNYloJ9Sqe616kKiBbcqLJKlbe6bJx8w8lKtX5Q86fkbQ+6Rrhago
sMcL8i8Dfl1VcEnnEbmWgaWd4s6w4T8495ukz0Wq0WWDb7Od/+AstAohvPexrcrBA83c0WMSxCHY
vf0Sc5BiCK9Q+r5I05LYtLCe+Q+vAG0/lF+KlMqWTd7mLLihb2e1k3Md65M0a3rwRkrjXTZGoyKM
OdLUYaPuSN5B/TAAn0Yy3I3G6B8VB8pAyafKWMcvkLNRGD7bEdOV7u+2BJo6bCkj5/NIms/55ubp
C3iL+yU6yQ8BSL3gOeC0Bqp7+jYWIloBhIGUJFu97lOCQfY5oTKxSRD35lTT7k/QfN7K0AkilYC0
719XvBdj6llaM8L3K7lme2M1vvcteJH978EaxcWPWj66L8nJ1MvYSlsnH3Y/I5ixYOtbDjlnk+Ta
0pv8wPyUAjE6k7tu27LHME1f9SCnP9xjBeC0bFP7pqENRr+rhL5VDmgHInqeLdfLO7cXyv12y8xo
U+bcqtiMCNUl9FbNvePtnaa7WRJ8X6cZLFSZaWy/CFFxI7EzPNaR4qoV26XMrQYOPXSachfVyFbx
mBG27q8u87v8roq4uAbHZDlqjRHO0J30pOGjIIDkmmNOEEtichZ/nOjq20eMVhUwoJTbjLyUcAet
Ha/P1PStPJBmnkXEKzwoPbdHEJO5YpzQg99PsHYejs+pD/Inn843WXA0NfaUOl3bNrudMi8SDAyC
O0EePlBC0FU3LGN5sUlKO9Qp54O/4l9uQzOA8g+irlXzdBgFlthiNsLiYCfgGQ1UzUMUlXy2A5R4
Rc649X8brvbowUYhWhA99icpeRNEpU8DeBxgPuMdig+5PYlAEwE/R9Z8G38Mg82fPbcEktUD0DaW
uYZrHJ4ppl+2Ybbk6eoTSx5fypH21ggMusqO3Cc18SL7mAqUhiuvfaoXWU1U4caxT8oa1bteC8Ew
Iwykqq8yMEoBFPbPfN0D1AoFsIrZOpFV0UQ+MvRQ7ETLpExGQRUiGiKb9iB+cAUAS2fr7srxeqeM
ZIPcF8Jkdiat6PdqPjS9nXSL2dCOG/ANk945VORrOgsMhO38sEGajQmej99Qu2VygsXCKzudzphM
oHmolLZUP1NT8Loj8aKfUtfLPiseBeLvxn7KgBwqvO/t1rCFQQRb+QhDnmmiZNKpr3/egw/6WSJd
0TEXPbDeGA2gueOAFdKVHU85XLft4JQ5iyQVAgSp1TaXNVviThJaQ+Ld78XJXeEP+/9rKuAqQ4/9
OiuMLnxgT5tNyzD6e2sSLEm0NpcNU3DRb4no/gZDfxW/AGTG13pqpJK1rz3kQo+HYBkEvYmggQG7
cJpaWxWfXgBlohknIylKhc3Qv1arWVj7fB2BkY/1OTyR6eoeEanAr/JF03xagXTy79aQ0/pTrV8Q
NKyKtmRQ5c1V2Pahq8tZ/KubYDy9DOUUWvxrqd/hUiKj9GswBlQ23P/JLnGavCu0zpcbViyJcPbO
cRxhz3ztStLtnntpjGtGuvrXh0h5u36lUWRV0B/4XsceAZAtZbyFCQch+aYS2+Z9/vlo/6QP3GrG
POdVmb7a2rJoc1/sVzgCgrZrO3+XMzT0zn6gS7DodcZ+E4TlBVfqciTd2OaLK99TnBriWJoket76
B5OrrGAJItcytQkAEdNXSeVpLXt3XxHQjDVR6Y4fSNPv3XXxOVsS8jwmJ6EbisjdAFs8wJdHRvuD
PZ1+it3gpg8ORaUEkRgqLWOd8SjkScqhO7UCOZbo+31IB3wDup+zAqP2jmhoc83k57+ieBMsT9HU
11TZU+fwp03oRiqHHz7IBkyM0MYTzgpsq5dT7f4whh/fzACB1NGUokI+3giMrbDKoiuuhtnv3LOv
RuRCrW6KSs62eFN+/MQE4uezQxrU4f7SzSwK+cPJ+PFPhr7XjI+eDBZ2JVi3jZ1jYI+U1ghmmvNp
MYA22vdp/yhxJWf7dq2i8VSi349EPJvCSZvixr43zltgmLxynqkV1tw5E2uUjTjTKddJBIwxiHHm
rcBNvyn+dUCw/CxYdmxaCzXDFya/Wb0AA95R+qbQRYa21BM8aIaOX6nhIYTWQurwc0sdwtmDEYmv
JMRYthKHK+jFF2Tk8kn/vW03ST+rfgsrh+ekAdwGcAP6HGt9D4R/NN0HiDDmy43f25BjDJWxV+M7
FL1Q83naBQrGkIln+8YV8DaSIPp2qyOeo4ulUykhMiz74cR6CDa7xKgfriRoMSyenoY7fTuCqVxu
UadLdRCryLX1Hzs6fT/sEi2sSipZRLMxTCimFWWsLAbZNlItjTZfHXvrUbFCsb2d7R7VxJdSf5WM
GFbzClpjxW+K4QdEoHUEhBV9Pc+L4XWeclh0C1rELw2R7zOgoELGsBvTO4rPS2UJQTHR8A+ESUSg
iHEae8RLiv3JVhZfO5noFxr9407jApxFxMbyMwrR4flJF0bDbbo2xG08Jd2ZfWJ+OVTH769/6KLo
EXr3m1IaRdg/HRuQOp+vrnBafiK0RItPrPrpD2weHN+hpUe/Kdq5dCh/1zLHbmwLJiFHK2NsHc/+
x3hxnw/hFGpgvf+kirPWU4fPDcWyOMxWG6lAfTCYZwxKXV76N4guPY72Vbth5k0rLFMmYfzHCE2+
143QyMxEqapqFoHWCx8vVj/DbK3x9sRRFVlw1kP87K5jt1qYZHqLpYR9qcxa1MFLvBTm/BgSwRvC
X7xgWUmvyJNM7RzNOmcP+7o3iqGix4XBKDgWAkEOjZuwEvAQPf1k2Tcj4uFBAuMRDR7OeE4mklZ6
Xpj2OfmuhvW37gv0VBD2pNyT49+FUkBLFcbvAD0y4MZ92/FiX8iL+rmX4y/CZXUuBecJuxOIys//
N2bCG3E59ofAMB6pyJbwThcGtsJpF2cP+wSwl8KKL1s46kyyKApd3vMrgyq7VZuVcHzMB82N9ce7
ojIygKWyZUha0RKM3/etSuI7QxBZRYKBXyjGqU5WWl+JG8w6G5Tli292ckrOd/zoH9A6YxoUHME7
nJaUAyRO6CHqq8Xu7PhWVbQcN3O7F69cgHzDm4bGLLW1gbOshxafn7o2YuJ+VcceyX9onWwxyozx
5YJXgTACa2JftBivf5qIPGBirz/vrxBD4+w4RySxJNs1H14t70OrU5hCVawXltohIGkscM+9qdFT
R34cUbkvOrjdsKr7dQblvEI6Ih3vZQOYItd9sCayY5uLOQXuWL0at4e4Ym3CbEoQ8vcCDPStm1Ps
GdAPtULIqW+PVUM5YmqsOO8JPxfMeQAZpTOWePIZbgdtS7st3aD57igRf7zJjWRMN7+txji53M7C
M/XAJmb77PApnV8sywlawRc8iZ4++0Dd8O3CzZ3/ykGsGh6DdqjcXZFWOmDWq9wM201rATbJMG1j
F4HkgyMv0QmRJgNO9f+UfABQtlx4ONYGAK7XyjzTKNRAREWKPgQePi0LcoghlyWv1MpDxdg8aFd1
iFX/Expv+/7FEN9VL/Zyg8iLAMD6vU0CvMgPNDy7XfZgM3vVQ4v+S7+9cgyBFBAwVoAvT1V9ZfOm
IdFRl09z+DbquvtIO5QK/Uc7pxPbWPN7NVsmQqDnTE4E/psa7xEy96/o11XsDUgXMfmT5+SdcRjf
nr/svcxCaDsc3it4IUZmu3Boy4GkIcmhotzGpdNCw5SsiDW5XF3dYef+H4MbNqTzfzq07l6XCl9t
KJWKYar/lsB2Rq3AXG8Wx0E35gNAEjwryKdV6qHPGrii84Sls9FwY5tIETkKluwZCS18zwSwrqyU
ejgILr6JXigwDIT3adb4mreY2P1+Kb4NsaVmyh25EuaqkM+F66Pl0mCAmCLhE5iXyCAUSUa2vtNN
cw8qpj86/HUSnsHUUCUMXgynyFZkP7tQqi+7rdm/9nCeiDOaIBkR5liX0g5zV9VJF9F5lvX58sIW
r9lIKtZZic2U8LSrry9/KgreyzRDGWZJGg9to8Q+M284iRuzdC6lFkQEvpSq9VqyeXmuhg6T4rHz
GnZTZ41QLYlc9/Q1K99/dFmP+m8dFKPHFRnzYd/UB8KhVybCvX22QzSFYn1CwnS9Z3UyXViV8Dyd
nQ8pNeJpcHkwKfrvseM2hXHAmBGRML8s0pXAPGJCuhxC7Qvo5lbLMKCu9KnsnsFDtL9YQO12ECkW
0KJiyFwy8m4oA1bm8/yszmtE50p2PKIa8liYHKotMxOnsXyBnnpz4dLGMJr0yPToJN/TU55rW9YN
ALMzvVoehniuPlaufcnhaYcco5vsqqJk9Yp+gSi4LA3KOOPrvhEyF0uKC7W3WYCYci5emtMzS75i
RrsaGV4XSNAjDTFkYG/zFw/+2Q1U95g0I8I9IO58PSAhqj2cDbvbHp5tTDnk6c+LV1fyC1r71FjL
LGD1CnbDYr/q2UfrGiD9YKHVZEZmOY97on+eZP58nu4ukII6BnRw3gRcfphHwNwzRbw67NI6cBqB
v9Y7+gLABGwro34a9Rc+QgHnqAg4Oe0KJH4SOO7ogx6YHoAuaoPj55xn4xR1UYTnU+m0BIRdKkBn
rUlic8Fh/XA21w==
`protect end_protected
