`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RkJCPNLzlO4rlRcNX8uuAF+Io1iRaXwBxe+olneBlwaDHLGxEGW6oqJxYb7rbVdOoU0Okesw0gzP
DWVNM6/MZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WPrVds5i9DeXqDq772sZHSJapzqNQWanz27I623kca7aWoQp51yj4JBJqsQmRz3mNNOE7IOKUgeZ
HWOQMD9wcojdLZQ8NH7ZDJCyC+piElkMFioqJ0WewjNTvBcyMSleVa8AOa0K2QmyntAdZPx4zdpU
OM03BSAZzn6JUt0xgA8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hKMYZEJhnoDdhjDVmPNpUYhZUKmJWI0StlvMjuR3yz6LWQ+NkJ1/R9uVlYDOum8J8oQXDSJonejh
wlxxUAA1oCgCzu4Ax7SlAFGhEF9RXaz6peuTInkTIoYoAJODcpnFTu2jljBbyEr7KCWc9KzlkUgK
lMFSw2+5y38MDW1az0c=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OJVfEhdN9pENxPVg/JJrel1mPAsKN7VMEXNGrgbFLGNDrfAApXU7nvDL1MwT4lZ/GP2iUgivjXmI
ABykOz2PHEbh/yuaHnUJI4QlblKIXdK/2IDxye2uo+YTLzCJuI6pIpTibT8WOfBccahIaEuhMopk
szKNbIz30A0oDIiGQWqknU/LeDuIb0zmUWU3Jq4jo/pO6RxNbDKlo1Yprz9iiHWhD3rlLIqzhQKQ
SlE9wiKdrKTo5ycMDmrGL+mj6CnMlqKtjZbt7m+LuV4PV3CSwA2hrHRsM89MO6SQPMzdDkjYndn9
Y82zcCS1PQjjhzel7jldyXEFxXT16l62eTZvuw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T6F7Gjg0JJAo/UfPkXZFzr4ELZ7l1SHeOGNb6WpuCbMK2KNxXpbRBFkSWTUEuIA1OKymhhZr17RG
tlhHunLdopY9rQgupi686lpZYnVC00TM6/1YiXomU81njIEiouDuHgpoHKjyskr3S21+aecsktAn
DtioiHZVVzCFqEV1ZaldHs5YB1Qnga8Zh6EreBtoU5Z8DUNxjcRK4V5MR5BFvQ6nR9vM4cApiqsH
8YbcpTe7pIMC10MHQsSxKJOLs2mmfMCV5mrlYacQTLdyrPa7i4r/8kIBnr7e+HqMTW5+gwqo292G
e2wi2IG2hPch+IuhFdTbNJiPF32UYrGcTzJGyQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PvK0sQp2fs0U2MjmxRkN76kEfRufpUAlc3PySszez8Q6pDzXOzsdmhhfnz06EgR2T13OilUUwXd0
sEGPgEuMjbj4Df54H0jiATYMJCIgLscMoiMYdZc5kXlzBGgYvN4ysYZnnblQyOgW6MTkS2pvjT5X
T7+O/rnWtW7R7twplp71O6aXqoI9bKvSk9jl4tQFTlJj6AWW6l3jeykszudHRwoAJEj5mkhjkDS8
9InEGmMwi2Le6MWKesPCPocf/KcZsvVpbCIUzKgr+jTEVcFR+aDSnwnpIz6eRa6LlWFzrrj3V+xJ
/cCF5uvchlLNlis+tZQdIpgOzPns4KhbvlaMyA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63104)
`protect data_block
mgnxztHCYq8mua+fEy1zdGyx0pyplZvNUWLvJGRpT+sfWs5NFOM0CCCaQFTi4duIXvU0hybxgZE2
gmfveVjAvHgERcTfprz2Hfhw3Ubun+SgK+tHoRrOP657nA/QzCdxkC4k2ZUC+Zqy29QY2j25kPtD
dJe4hVyNa1yVbEfdj7u+ZPxCVzfg4u3ypa6h5yb2LAFzfywHat1waRr2DTXCUeMCGLI1m956hqD0
DqxJ6Pc8CXz6VqJVUvRdH9Rp2bTd7mbrRl4pt1CeNM8ej0wdBhfvs2bsxv/m5ivuLS1lp5nf0ufo
9XInFE6OkZyVpIZ/xx0gRgrIyaBbAqNTIph+/HjCqoldcHx63Fyt+PHLEol930zcLL5va0sJ2aXd
l2eCptbtmHj+DQxxbtlOOoh+oRj91HV80phQicOiA1QXsyPrudc+Qtym0SZCRnrWe6CdqJSNsLZ/
f69g15IjvRApDw0ldW1bjt/s7X2Ay/ewzaNKFgRKkRD9DzCeE5qHJAv8I4F4dYTXA3bUami0rBZO
qedcVERuVONT5f4AncCV+ILhj8jMqOjBz1uRnzbw1rKZRYcjfh6wAGzBlrOfS+0Xp1FEZaCQbfrg
jvu7BIsE8Gp//keNCIV+jF4aiFlYtxOkKat8h4GLm2UTWkcRbufyqLzIyefH7PK7gm4AUL48fX2I
IyePe/zHk9k1o6/Smbsbx3ctCQCdN7zs5qVD22S5QMmBiv/YsGH1JcNKSAks+a7Q0AYxdXaHLQhS
AjO7bn4pkBZAuuxJRSzddp4/0Omp7g9wTAH1UfuqIoUMvV8jwVyW5iidHN0AcmRsw3XzXM9ppJf6
KXdGBE8AWRi3wcx3kvuiN+m4dL7y1CLz4RUl+b/uzAmw1DUcwlq4sAhrNdUe3BNhY0i8psded938
fCOuecxD7Nx1tsQEujt/zMlr7bwyZVBc4p+HdU7jLlVMkXCqB1xSjxIyad+arn0OW212A/IvtR7U
zO+nzF7dTgJRDcYzGWaDn/mOpvOWH0TIS7Ia9lo15uNCe3i/z1EP2yvR+vUz9warvQW8dA12QSYD
GbzRpeWOO9anBePPeaAeh1tjJRW6pp7PQB6AoIUznUBnkgMAp+RxHOsRRM5GedT/IliW8wXps3Ma
ZweLFpz3wTMwxf/KEAe/pmTZa2uGK5QbIudP9IFJ1thhHwF8M44ItPf56YwmeVWODMHhr/PPqKyh
q9AAQvQ+v5RdRKpIZjrduFK0WwTV8OCKJi+BbNmWdSvQvCrCDtqMBeGLmSN1WPfU8QlmGWKL9DzV
z6yzH7PbgPvyqJ6NNChpT4Jm9RHK+7854Hl2hOFIfHD84zRuoGLkfvrB+R9WEplZr7XlgrIoCS2/
l/FUR0nNX5DzXadVY2GlBwtfsUojIG7x2vl+k9n9XsZK9JYyyCAp+bYsjOXbtHt82u1zK9eGtpFM
a+AGEe4eW0eGvE5Egy/wb0p2XFB3Ay6IE27eiPvk2lMP954fdI/2TiVlSD0FQp+I/k9WQCliY3Dj
1OaBWLhKareT6TaYxxqNByZeWGNA9Kc92TkuujpUorqTBKSDRegMaV8xufOSZvphMDsCp6i8BqNV
VfZhwEeX27mAykkzIg8rP9GNBicCAMw+FwZ5lqLlgKGMnPq9dYUrmN/2CumP12+CvpAl4R2y9dIP
IuFBcY8FUy9OalELo4WihNIpkBKOBlsVpqZ3mDddEfsLY3muO/Lh94l9dVd7OZlIhIzW2OCqc5nN
Tk9sfxSAsT90LUqDRiDh7OdDk9wI9NxDG3CiS5r9Savr2Xg4jfDe80y5Bgjjb3oHFDG+cUk+H6f3
Ui4Zl9ZfVsem78iJ/bjYTQivO0d776KmJzq4paM3c1PVhYopiUFFkw26dhcvrepFOB1kJs3eP3Zg
8/GiXuaJCvH7lt0ey1pw3CgfcWm5JgYqZL7viWKFP0H+DG28FfKfap5w9wvsWMDD7eO75LYkniW6
ICl5hXG4UDChDYOAsJsohvnxHidTy5CXLo2AreKKp5A3wYiF6o7e5BwZXZj+XrqhrBDJkkKBX2Wo
7OOzqEY0yH2yXj/CpUkGAD8IQkgXZrktNlv0mk20YxdXUUjr05ZhCzwZ/2yhQynpSHmr4AP5zNdM
+oR2sjGfvZrhdegm2u3oh88Vk3GLOV9bNPwBAK4oULzouZEeKKCo7lCgEErYOcqbI/Qp1j4e3u5h
87JZl00SUm6OTFbnyaP/OxQPY3tfsiybyyWOpSgl+xAQRxidpD4+1N94pzDmBvN93UEkmCewhOoT
NFukBtpYxpskrZebV/8GjC4vQ+K0MO91q68ZGvDz1m2A4dPvJJly0A3CpK6JF4OQ5KPHcS6OuaKt
vo1TFLnGqx4Et+Nys6ZRLWvvojNlQE888uAinPZ9BDKqRBzk3VFUaBfaHrBEAhL7/IzV6iXb+Ssd
gwo3Hhhs1w7akygkLoldla19c6hG8A7T7ND4oDqws/x55uNzNf24RXdf1lacY1XaB4CZGjKv528Z
RCLEj2SUhXlDu/k+DGvF6mrSfbgcxX3Fp09IuXDV8mfAL5Ka++mHj2SXdxeP9wguiTRypR90mC7z
Dbib5UAzBI5HMFx9XGA9CjL5vhYogIbdlCa4jKmUUnSob9enMnn/N8oxMS6eF+gpO7qLcgYCnFy3
VL0bAqh6a0AwPB7CO9skoIgaEf436jWyemkJcOL12fgImcbL3lJhS67SVe7fVDJrb5SEAU7o2saS
82L4+uLrrO2V0udpxkP9qc+9FVSiyX+noUpEzIsTu/Xr6yc0g/IBs0Okzwnio5ekbYJ5CDyR9szs
YQbmiaO2Xhv7O9XeshczgXYDu975dV6DvjYJTKFPT76B0+iXJmjE9CPfQ9SkyugyaV5RWzELiIrO
CVtLP9ssKcFlVA/Oz54qxdgh6+myppIrwkmeoBnXAN9t1E82Msc4hZD/lGLIJggeqdux+Z4xAzVY
wP5rQiRLrWLlbQh0sIyFI0rgLdus4FqEve8skWLUn+JPLEIIsxHeUD5SB3eF8U3sJ8NtPVGjW15T
qw07aEjMz9faoAmbOFjfCEzemQwrOAOfeQjn48uYSTm1iYzRLFaj4rYwarMuZXddlYtdci9UTPh4
S26pjarUERqVMjupBp3bidqVNTtgGiaHEf8CMglGwNxgh0fE7FqoZ7rdCqKiUcEYtqPyOUKbKwEN
6ZYdH6+v3KiNg5APN9tYVrx+isPYcfDsxyzE5dgOD7bB7FAgEFGuIzLsEvNtppbXFfHfSk9teXuk
b6B3kaI1Zp87wywmhSWJEeX+qTJhjf1SjdAcdjVAc0ENUcgOnXWPAvX534kXCEJv8q2I7soc1pM7
0lwjH+zrop1xBrOvZihZ1mh6U8TcH3d8uFItxiX3MQ5H4JkVdiZPHqFipD39Bc1vcc1foSmvkTiS
wwesh2MwSazBaymG7P6mRr9Uk0umzlqh3VcI4+zerXXJG1sMNjT8PYIMtLnMVcoWH0eU4KJK+KIW
fL7tTuIg2FWFU70BY9PvPiwQ8NwFM3DYWTE8HOqfxGZlDku9Eh1lY2KfWql7T15B2IsCqI75cc0N
5LqFHx86xeu5BmKPYX5j9PqUt31yhsdrW9uFF6OYI16Rj6TquttKlHdLMW5haeE49a4F2khQUq/B
IXEWjYQGpRgguUJ1ydhbfne5q8p34p6sBOpf+PNK7i3PrZvHVAQ7s+wFUcWm11bg3b+KI936HahA
u/rGKyqRBdX0KPyK1Oc37Ou4X/jwdthUI9aPIUbRJgIDbCOFvmsALuqtHCm1Wt9bdSGanSUgwZNc
ex78lhXkDqsCQEqPEp21/M2ORECji6zG6TOf8ol1gZmdAwEtFqHL7B8tqYpvB1rWdxYCiIPfpTbN
S1W7cUmDG2bGuT8RyCxDM5giqKVtSlkzQVwOaEvnsWCIHzcH5nqeyg/PnT4PrGsEhs+3jpVF+GaH
uQ7BVZqie59PTv0O7QmQgc9vlJ5sFgdKFF9rPa6qzad/u3Lsfw14i30gBEfLjheG5t0Yl72YgMLZ
owgUKEjX1lq2zYFQrDp8eZH5PknONWKv54n2+jfb8MbCCUWPHnmOXkMLuXeE2iPYXjmZwqLvO3Du
fglKJC+hIMYnFoqVjdAhMwOz3j0i8lWJQ4XOXbqQqNl7XoA1sYvsC6rmHUi3Syh/oyzHlYO7TkiK
+nGT/rbo8CeyZW3hcvfTlT4TzQtIUaCtpoCM53uxmSZD/y6XW26tPgMqK9z4JkK60TrxdxIvV+qX
hXWb7I/HF88yGCqfGeFxvMLRUqfqHzmdyOA7KS1vjKZPwBEeyjB8mm/GcpNZV25H79ueKcMCPoFJ
WQGIvyPFISA40fZ0g2SxyAKAyKVZpJKQxXjmFPTKDlM6c3xN/N6bGmI+uSPBL0Em+n+h6l9P06Gt
k1Yin8JLh50i+ciAzCJhbMWbWtwFNTHaxC5hXNRSnDHqqnC4gJSXhmdAZKOfQz89DVR7WQweOStK
kg8hM/PlTqsgHEIRxyn8ftNvp0mTssWlnFF9qPf6KcRVzFcw9POmo05uM4HwOg/RiuUBUXscsc7I
63w3RnJVADDr+OlRiMuGLQf2zkM6XIba7MaxIgVFJqom4UWSuKQP2KRE9CNjjFuFdkiH7+3VCvwE
s1xMcSi+efvQ+SzpxeXMX9uU2nebKo4ZmZan12ZHBCLWMhqZvC5i3jNJGvCS2LEcounA+sPXpvZP
FcY3I+WqzU1Vb8I8Rt8m5AAHLbCysyw0P4umJk+ZyjYQ4FL2L7VtsJt99FW5U+PlD6eOgDaPG/Uo
UbvS8HfUdAd1TWItMUH7B9qXzq9pwZHKEB7fkQosmYcj1EXDUIbfkXeR/cg9HeimOceiTNuCC0tq
+ZUvvaPDHwdHeMyl3OmJUxtViKFFwUeNk7mUU8PF4imryYNK/y7bqsv1fuMmljncLTKu2FsTsg4b
rNiFbPQPfEg+czkE46BOu2yYeAAXR3NtRj8sL7ZHaPkvZ//qanTWBRFJ8PaStDR0e3GRNo3xc76u
y33fnSWGWqGqxMhD1w8BfoiLbKNoPE1Q5PLxRUKvUtCCo8zzY1QIYLFG94p7ymdEJDkL7KUml15k
aatrS0mcFJozYtQg1APnRiAz7UmSLA1PgA1HFo/5xhWY8JxJOD35aSbAsk6aso3f0+rlhzbahTPN
Ygvyqa2PGM50LufGAuiEJtp42JJ5N/HnLBMXTpc3XLllnuDzH3drCGmQvvLoWa3GXw3zfSX88ws6
SsY655b3XvGL7bY0kpAexBzwyBQHVZnCLmL8D0tk3FSJL8W09C4unI4QqUv4sCOYO30MKNfmlxMl
wx/6PUn43KurAJ4jdZK8Fpfb46PE+DAh3PFX6/l3MCQ/xafvTDG8+/ZksuYnKy7Kb717armyeaBJ
6CIxkxFGZ5Yi7ruzwQFifVZYt2JFLeJFpHOQH9zxMnvTdTi7f+TLhP2VZWIpweFtEP44NcKyNB2Q
OmPi2J6EOEaTfxAZb650nwb866D8xymTANOjHnrM3pzixPDtggEYXOErVIsD3h70WyjVTCxMPEiJ
iGNrA9XcwXgIy1Hu+bG+ll9tgHZyGDFr5YltJI7VK4CYc8u8lSK3XLlf7qTT8qU0XU1XZDJejzUI
kGiLTaaipOTNoJdUBNORS/6kI1wR9VKMrJt05KFOzo1ayPVDVJ8DOJKVHrRsXWtW4OcIRlBZLAdl
2oeUzgBJ1piCVgmFyQ2g/+XXBBJ5MdaLT9WZXI/l1P5vwbY/HNb+EjLA8++AXL2ZraNFqydLp3zY
d2TObF4leMYu4yykshOuQGHap6AiNEJGQgRK2dY3gkIksFWGJsLpaasXcEoz4IhxmZsuLXneWwRY
y0naMcKc+OSDTuytANRhrxGIhPLbWauuQClquienWfvp8m/6CmxFH4itHGKOqc1id1lPMc6CyM3i
36HL2/mkCq1cCHrJgwK04h8vrl5q6dYAr2d5JPGYN5kCUuZpABs22HF6GwS8CdMGuI99Xz+K0jCa
BByBxLpNpZcu0ucZXZRTyjeAr4R658qJZp3ClHhbIChyIMUhFGGZFS/06Ojdz2gSXAAIk+07lHMx
wbi0ter0/9y99zGYtXgwcFUVyowuk5/6UVZNUb3JfEn1gD9peVNDgDHGmnc84bID9Wg3O00Dw3TN
GM2o7J6hLLZ4jx5SMvRUIRylAW1VS2rFksZym1sNbloHto1peosnuLqrxSX3fCLEhInDHgGmAlDt
xB9pR9dCauPtH8CHLJRepORizzvDZmQWybC4JzhJYuSTbyoMXl86oZgbTpxIWYPJ/9/0l4zRqNd9
PEKnO5WJJse5Xhw4nf7fFdkITnYSjsZwio7uSrCMagsErqOdjeKdPz0S9ljpNm0t4M73El70tn4z
3iWMSQFbsXDcJQy2vvopg+nu8OsYrM4YiuyqnF9lsniJxD2SKBC/mkY4PwMUJl9SDd0O8hofOExG
sTErjQvmbRdtG9aGmbamqZDxMHdkCRjfKHBK6F3RFIqtdl48IUOrq9J0wVdnumRe083mltYQPEBW
6sJvfPqqzL3M7Y7qd6xsRpfAEB4hsdUHH2dLc7yOzZXeEkC9iZvMG0DHjLaWEhM57Lq1dcv0tqj+
z76dZL/QD9wIuVpH4OO3IRlx+ituA7UuuitzruJ3J0xwLiHZ7O8aiEkDMuIEpso0cK+jMGmX4v4P
KdcFHx0n7ytcSyIWBUsD9auLrSdOYi+cE5LMgXbqXk7GxPup6zwT0PzzZCjHjqyN1uqS+tc0Tc9t
s+yDy906J9UKJREdkk/nbv/XJWkPjMtsWzmLZazjgprOshRiYEAoy1/WtwLv3qAW5O2OVMdunvha
g3Bdbr6ERlWd6bf3RAPBJevOb7OGHSlza53Z14mCP/ZzGEPm0nmp+iaVObTxsEZ9RVXqAvDbcsIe
HGw78S9cATVQefuXmCSevU4qVDBpzUhD9B+i4lmWXfdIk4VCfxl57mStHsHbH5ZEvpAknjCZK05K
t68/BiV0Etrb/HStq7urLsr8ZKxcTqXwhaHr7735jP6pYJK6LkJ7IFKJKBKpVe1YO0Lm8QYqlr7+
TWMs/VeQgmbydE8VXNEpAA6VWZqaLguKRb7ZhzkKkxq/U5sIF7CIpYdzMog7dKIu3v7zq14gWrO0
o1XybFqAo3mrtAlqv23ACyjxWna53XiZ4P2+tOH3gwImJaf9v9a368ld93zkb8321ZQAi7rRi8wm
vbKvBmRKrHgmKaPwnhmstRrI318S2ykWaCkbx3cfUc425KyZkBElmgHVvKIqY0/3ewYsRTgMMLZ7
fNXWrdsnywwXWpdTg5xJxyUhZHjrmaMjybOIsIkTv5B5fJOwZB2caoruL1u/ReZL0suhGfWVhcx7
cx0+5advgUyyN/Wsu5F4FbVrI6c13ZY4QxtWkZPY9m4v0G/sijBy6ZeoxeqfI8xv8Dd+A3vHm6yt
LH5JPc5F7MHDMHjtuskB7sQdNaOEMSpacr7N+SQe+ZRoto4X8MpSsNVOqrdle+C2Q3WueK8fl4Cn
pIWWSiZVdFMAF52QN8f0JgaZMnLgDkgBU6rYbKLsqjFJWuzw1z8Kcm3HFU+IlZWj7WormVTh4MqH
ro2FWtJSyE46hP6G8XpWy6DTud3IotA1Qgl7zILXB/HUaEUN33VtW90t5cEb7Ys5YN5zNVFtHblU
168o343zrOfP9bq+y1ppIMjnFc7s8/1jP/AZwLkJUOtPwf10dvB7sJe91MjI8Ot+ItrQBru9ZBS9
bJ3IFhmphN71Tope7QGx6U9yqvEy8TJHz/MSsi0wJS/lDNXe+xBIiS8Xv0QlKBM/sJbQhMTrKZXS
b0i9B8eP9CR5paA8oI/LM+xJAiFqn7JXkt8QslC8/FqsZm/+G+LJNxOEV0iq813PB2bxIMtdJog2
K6h/VhXHnEXH37yQYuZCPbDZftT/BJykQHd6pI63l09/K/nxVCbBwIAPFJwH6wcSTpMjEjhMmO3f
LmMEvWdxWb+1120xFv3zVTDM5vsQN4IlVHTOZxQyJCe0JyHC2LV21eNb6sVhBQJBwC4jMHGJoFEJ
LoTPmvvdI7kArKuRk52yjI2TPRU4t0dblD8xE0ao3GQmYbUIpPwCy5lpfxzIRsC0lcn0lyTw4tnB
fTD/Ski685yoNeQDsiLGJdXFkkD5oVMCOuZLKCIlZ4pOLUiBTgyaNTiWu1E0wMCapMVGQgqfCTyg
rnRFpCTPcmdRD5+bn6lLTWaoBACrgOEdf7bi4toDhWzyyhtGszlmo5MLzluO/t0WIxsa5svbcQqs
epYyEgN9XjRz5X1rqygRzXrivjXNzUtgFIZxBl9SOzKVGh1fuEDE9EfMvepMrbJPo7U4FM6VscuF
dQRXvgRolIKf2SJ45yjq8Rcq+wfTQ9ekwQrZjDoiZJ8T8eLH1xKGtT1HNcmQNTQZAYdp8gnsi08W
etiNAazQJPlGHmjVyu/2XOUT/bM9F0ppzlP0onbj+M/58pPtK7yVD7AYC4oDZYluhzm++GnYPKMT
vTnkuDtp3u+d2tllOG2MaL23Ybs0YtQ93p78L9wgOMk8txFeM2eCu5Eba0EbwOejt63lPUdmjAWM
mPQRDLY+x/WnU8id1GWxb8gfkMjSp/A8aJVnH91Ao1DZs0XWFZiyRQYpQNwO/1EFOw/tn4WhXblK
Dl/kkqzzveXB0FA3EOrKxN5bS923TkgDVtfZpl+lGAWTMM6Gff0CMTBQwxss2b4+P63h84lN5hPV
+RdOBrfB7W23irOhWqktPD1Zg6IEtiXofuhKfuIOWHIKzYj+vPlwijJ8cY9GrLEGLv7/U87Fq7Qw
Ga64G/tG4FBIhkp0lJsGPdcoFHbvdj/TQlCAPdFic1G8SQx3jfmy7XcFH+b/HY4Odc03JIhjgUWC
26rCFwBAwoiO23MApGXSY/RLklCqw4CBDb869lH0i0gTISk8DGWETZvJwAauHeG4MCguCErXQSaS
pctHFDUQ2OBQBJ5uX6c9nUhvLYtNeSCJZzVDjbxfQUvCONYW0jI4xvAQfwrWlrBDYTnrj8Ud3fl4
ATa1YVL1Fhscs/Jr4PtFUpszFYKT+rdloLi1P9WWI0wVwsBein9xMByy6QIISoDRO6DMF9RdNWMa
jUyquWmGU9RKLFtsCquVrWswDAeFGP3LtzWbMh5jI5wNCoAAFZ7GAbOV1gHPQowdnHAcYCGVfphx
RjnT2mcoZ3LfIXL1g9W/JBEZBIulhKj9TH6JMku1F1DAGFMDJSLf1Mg45fkb0Q10uwrVQFsE6TdQ
9FAFI2Lbrz8jQwSVUexBjGoZqv1Jii0YW0vt51nniu88S7YVZaGe0lJMwE+sr1xDP9mrtBwqVOm9
uK6dnGflP3+w2h8u2xbsrb1CjaPr2VAcC10b4oAg0V52npAC5wtJuZChI9DciTDQIw9crR0xgOnk
ZnwIRxQkcinU8HpFfpbNi7MDWND3jqGQz/S0J8YVkUH3V0TVIoLuOv6YMrJ2UZwrehyRNpVc+6WF
5MZekp53KnH4GpMWc0XbvBHDrmejSWqMiZv9uB51pjA0Z/UsSVSnkE0yODZ9D/1JudpvhpvAqaRW
r4WGuIOHLcDKTr1ljk6f6mXHT2FO+E4QtspFa/OGhJzATrESxOZwhOnNYkFPAjRQmgq9L+p2k8at
UVzAMFUKX/ZJliukgTWDK98cSFubqzVb8RDy1iYM7iJBqwx7KUDg+sm75tBNFYWWBof38tacQfhE
MtcJWuPF0wwKvgudt/qx5JJURDtZUYz4oHQCaIhE/wFHk5ocQvCC7m1SUujFKa7JkBk8xiGheb0J
tSvLATQVrOXImrH/Qqjc9GSlIYEOp1yVwqib5wjXK+ouqcda6qRRI2QqFqKDS6iQtqhUot9EnacH
wTnEr45xj/fEpVFwUgYtXQR8UhwTuMCyRLger5kJ6W27icA98nE7Q0x+s/a+UnW6PUo3l6lvan9x
bwW8nS/kPz2MLTQysl1SgYu98hx+KzkyYBIj30dGY451+4Zn7aPZ14WSaPt09cm1HgslEFrHaEym
PdDLYYVO/r8nf7dIFq2qOTmIkKi1a828eJo65i1GnTUsXlbDrfKkYK8o0dq92IaEWlKKKBn+444H
0pkvNP4PZlPz9A1ngyr99AplBuYKntHZdLK/rhqqKO1DCiOU7tMwi/t5WdwH8TdKg1K/Q/j3wrps
E+npT4sTXKlLVHeiPuq7ggvJqnyuckBxc8HTHti2iXLRm+cwmBMg9CTjtaAaJwY0g4V4rN3Y+q1T
p1CIDVSW35jviKOftFEu7mqhas5URBWrWTTsfFWnFaARhXX66wLtKMq9xk5LUw8OgP3mAstyGswi
WYWjFgIdl2sR39vSzbk29azkD8cz1/YFbF9+HrzAaoKJcQPfoWBe58s0a1yRtYQlf5j7RFSWpY9t
+i85yD1Jjwh3zSlNbB3+7GR604Nd9nYfB31o1/xg6zDDl1kViDu5jnbn6aUmzKpoJpeyXBdG6ONj
lGSlUN4G2XiquLxOnzaluNTmRrOkyDroNWrlxZhiAYB2jbce0SXAoWOYUqhtuDy8ZES2aFqKAYur
C4eWR6BxFCWcI85EQ3SiqofGLgusI6/UiJkPf4JW6EbJGAoyQSQ2BEWmzdZk0Y/wTiOwyiktlIxT
Zku70llbmux7IJaYkOjiZgFTnnTS9787BHhsayCMRwd4MDQLjXfOGnSEYPL4XL6XKhGy6Ydynb2T
fk0ywI9684HU0hvVYxcsv0kRMh9Uu7ZS8bt9tngUWdnOZEZz/QrgE+lJCrLsj8o6u6DMOVfE2nRG
slqir4yJeUkk7zg9dQE6xBtycUnC1TCB1CLSYrc0DhFcNasLIIq45pnJFnPixFl/HM6e3motdLEG
LQVKREAIpokTPj1eQeZS5wJv/SpViInT9ms+ORZuH8ubOgLrSGZ2ZE/vAiSyLcimzg0IZslXDS7I
/HoQfmyewKOx3WVbG8+7iyDFzu5lNgeWT7E23PT2WrPqTb5nXguDPDhLyolgXwSDXf2DWwrvP3Tr
5uNKw+PePbaYWDAJqqkHIa2pf/w4wfK4XuUE76CnUXoU0MBl1gYfWnWJ385MfsWvX9hVGxxcnj1P
hUwOfd7WeBaFH0SeKAswzX+wUgwxZJ/hiIa00tUyoEiFjdKykzDHwGtI0mf/GgMCBXt3xEBk9yTk
2pOF97Eo/ejLfBCvwnAtX8dS++HeAa48yWWvYMbamKt53QrjAC2qBC+xC3+S/8pt54vzLmKWk/gh
xXDIpmidAw/wR/AyMuAFEBoPTWR3BZMYfyDvPDTS882oJeNLkgeWZLgdUzxcNbVXIzm5xRXgPZu+
s9zKUXM9C3aubZZEh+vqjO5k4rSj4bvGo9RflmfEA95I3AgoJdL3cXtg1at5xWPYY2C68n7XhWEZ
AHT7YQkM65tao2Ch+SzH+gQwVv6s90IbNL5KmxxxyDfO79eqSwxa+Wtw/s3unpgP+AEh3SKkb/qg
AL2G9rbP4vfSW1eStESaMDE4W1BZ0cIrNsABbo7+W98i98QX4BwuCR1LfMjqEV+wpsbBn/Ko0Y12
S++UGMDc3vgQeW3kpFj4X4Lfig3MntWkiEO31tOrb7UJoPAmn2KOOhzidZ8k2LCpUWH73OWXjQzb
tw8FA23F2Q8S0ahAXqa4QkNupTnTbrHDACNkOe9tp/hrgfr4M8IzrwOHuOG1RVLu1PbK4aJIQ87U
Q04T7sekTdUdpWYyJ01Kxyqfq9GtvYAH/0/poIgwUt3fOMiR4NrjkLVESlxrsUcIuCs6esf8BJqA
dkXdZtvp9bbtaEnTDlGCIKS7fyoYhxGO0hOF1MSOYckTNCU7bUscZ8fzH1Tm9N54fDWnIh8kce2o
33RP7+8L/y7LJaMZu90Afad/MQfzn+eZvQw11WRzRYpzI54wQEPDbCb6zNDrFTOpyuTkTHb6ZLoc
oDe2jzWw2wrm70JVC2FVhRK1IE3DCXVKAhrUi1UUblZJgpLw7B3pLQlicb8pQBS61C38PJUuOEEY
ymEIZ7ozG9TqeVNQEG74jylSCLMPZUIk4A0EjI4hVSxBOrK4Lj7ds62UDteNOX5JqZfIvhAsA/3W
mFcB3DLdlKhP5/d7UKcEdHGV6GUtonHtGs0gsm7zPbVr7mqiUMHJMYQbCqr8JQna4Xr30c+wnPR/
I3AXlCFCqzge9hvhtIwd3I2NYHVlSVQXFmMRt1JU9XBcaNpydW5+ksJCTJ4AUHKR3oVTdP6QWsa8
kfstvDG+o8rlnQSK4WBbVy+Xvatq9jtZwhXVqiInuSljM4Xd3n7Uur0L1Iwww5UT6OUx/8wwiTqC
Wye6hD3X4rghUAMKT2HJBxz5XJml37jj+UW1lI05oJFGRpz0fnrqkGYv+PKFj686mJeHa1vYSWag
d9MmFfmlpJUJv5mp91t1wbrgZ7tyPcAPNHaNA3cKHjtcWU8JWFik9vcR3PPwblsbaNtfpmFj8eTU
5uP0/g1UYN9xCqxUgApL3uEM7NGUCBTYtFyReCwycSXTEbiGVislGj49W3YbvKWypmISpVFsVc1L
UcUQ8bDo4i7x6UvjXJHMNocZX/f6MjE87DvE/nDyoEaXM8cOnMYimYBOZi5Eya1WqQHFelRdN1Qr
ADeNoF9IyidbZkxiGR6dO/usMGD3Z3L0xOH8SudBh2D0zN7FYhQc1bgipuy5zMsMi8v4zGYNXjAV
FbWei2SdBoSYNSLHs4xX3VZv9hkv1YlDpRVdPgskggau/AFW1Zy2X4JWrFL1JjlGAtD5jt+i6jU/
qbH1s2DPMNtqu4Pedl2LcGyM1ef1MkGKhhkSSG6E+2ZjEdVpxSuBGcu4nqy/bkynn7AkJTCw6SyI
VOkyy7GlG7oOMLqrjHoo4TzESagWnY88CBzpkchkgrRd2ZelIpaXOTMLIDfGzjg6wA+giHLjqqPG
tRe5HZ8ohSbKt712gFraAjKXR4U3Zk3vHvu3Y913zomNixRwozlkB26vbnrxd5xg7zfF1DdgfaqU
ssd8PyOJmQ8KyWQ9JkyJT5J6N/Eo6mNBaGn01cEDcnkEFcpQO+speWLCRCObPLrrqhPNrYm+ZFHR
yrXr30Rs/oQQ6DtZ42zduQGCalGUCe205HBDCMtW56/YPDwfzBWkupY+J6Z/ZmWD9gAOncZXWs+W
cvdnrJhXGpQya5r80OLuZshN38XXx+5gsJ4mBXrM/vOz8KkLWVzqSDFgpG4Ok8b/ISRVSnulKMcp
At1zhJwjLrBOe3xBeiB2svc/7NZIj5vyo3cVeklWHvHyxX7L/P91iW0cjxD7fo8zJhEZEWvsoDlw
W32iS39oIjXcqC9JCZsO2Z1FF6iCXbTLKrRDoAwUrQqtaDNo4Hx79lB9lXTVUz36ghbSask+hoof
EPCMw3jsb41BloQxd9T0Iz2tSv6ROZYsS73KSmVm8J5zKoNxjZoi4T6gj2mgNR8pPck6RULDtYqZ
LOXk0CE+asvdkGX2YKX++0kNmO83LYispj43xaNf3acPdoFUL0OpK60JRM94Xq+22f3i41TVQCiX
l0Z5f81OfbMRGayEVcUbQXl4SGzLkGVF7DlkZ/ANFnh1eRw7VIdTvHnQB9WVZXo1nTuzXmjESvgB
mU3HZj0SA16bl4D++UsBb9KaOb2AfySglZOUhKhH7PCyJ+qgFg0j0LwQd8neeXHQkctQip7ij/NZ
fSnFsdzaLI29+3rAZh4yEUBTK0vp5rU2HMf206I8yTY1kiKqvVzvzkgkTc2fY+bXqfnU+x8JI1a/
XvRFOk+Q0Qj1zCrYB6N/lsx5kiqOnAiOe+Z4mgqneP27N4bnHveK2PyDa4TxWLVDG9F0w4Xr24Gm
nk9DowiiSecICPzjgUXMi/IY+lAOeprUuME4QR2QieXRnZEgv1b4ZNpIfe85rpESWaQTR1yXjrDK
86osG+XnelpSqHSqxc8hPMdSKh3PNH+/VKmOjUN8l9WoKR3ije0Oz8va0VltfzqtIhvARPrRNsEh
rxbMPg/fRpWjBmuU4On51OdF44Kk5DiRjp9P6IxMBNRcTehfMbhRSM75wS6YVGKH65Aloynip+DL
JnshFrMZlnxA556OuEsTqUhKCxfxuDk7gWMoRXJMQ83efZydcAKX2GiZ6uHfVkeqJqonPCEzQgAv
jpqVj1Cyvcx2GRf+JSeFY4OOfH6WTJxxxlXBEVOmzHGRDZCtcQSCyNNFGYhINOpxJMHK66ERVuc3
e27uPt541CGtsRxxkArpeRetrpC9EN1wuejibN8O5t6mBFlw+g6Bp+mb2co0SQuBVHFQz4gqPHYM
qqaOb8ur6xT9qAeh0bQeOJDt6QQ71HISEKH+r4UX5pe2llA3Z2iLROucIV0SdSokIarDFiKYLbJY
/wyOqDgmG5k3BKff2/c5mgVWhO+QyNMIXEk+0kwtJkAkZloiLOEifgVPlb7dYG4E3OtVGURI+JNq
XN5GAf/2EFdf3ubbzYS1I//3D5Hf0VHV2omyx9qsNNkgY0vQVwA2KrtcD1WiTi1q+6UFJr3F5bL/
bpdSpQvmNwaOwPqPTacKsWGm4AIy6b1eywvr01o58DmLc0AQmcSh7EUy+q2vlij/Y0A8Wy4oL1nk
4NCQSqzBCeetZtAfeUWpX1x+qVIaVvbvRndk1pnf+phQV6+m7ZxPxJ4dIyQEsIC6CkLPGNP4c3Iw
qAylA012V8IAytp4wBbe33kTxZx2GrPTv49VP4fO8C4meF0AjjZLdPCGFgTeJv+BK3P2UQm95Kh8
3AI96F4EMpKLe8mKqeKszOLKa1jVh38VjujtlUSWOG5tab1Y3yvYylA5f5GaVreJvz8KQeAyhOus
I/eyc+DBEHRL4VyzU11zcbTvZJrY+/CFx9uXmMuMeTPP8iBgLvxsjSWr78SKzFp6LmJcz4PG+CG7
NpfnDNjHmZHDxfrlgecM7lhJsrB6jVQFj0d+i0/AMa4/3Gh+yUrJaLczVM9Fp+i0hRgdz6BfoPLU
zp4/IeISBdJnVHhH2OjZR/ivWk2lxL+qo9YkP08a6H7qNsii4h9ZStIDJEXWaDqkhReyg3UJnHCa
PFljeASaH/S0j0LUVywC/eXC6YCLuDzX3dufxD9pMI/CRsEw4yzzk1iVqKvPCWzjKSQXd4wri5fv
2GDhDV25iArnTsfjildA2Y7LT5Fy4gUPRu+2P4HM5VXUjKkJg6B8uYQA2DtWg+TxSGR2FC3eZF/4
pkV6ZokfX3PMGT1Lh0IaKynIot6Z4AfagbkID9EFnM1/+by7U71FpCaUa/JlRXoH2OXdMLiV95jk
vn8jIamFtzjqIXt5KG1yMKmtwJ9fwpoSEiFLWtlK+nsPpt6fFTHm6v2KFvj8vxYNA3ucy/H5pYPL
rXKI/4NoBUOaJtZXc5njsFJ2oS/TliIwoYKn+MgZP5b4pSE4oACRynSNM+Od1Oknf+hnpY9m5+RK
/m0lLS5dOD3T5K3IeKKr5td6l9VaXyZa7wshXav4DyShNLbwZlDRnIQuh9IaQ2/KYdJnOEPPG+Vm
ZHM5VM/OAg99svUXWT+2KO03o9dXXlFcLwUP+JohJQ1YpY68bbp6nqa6IGF+HNNXu4rboeoVPXEM
nXBMfmJ+y21yp/AzXNulV8c78VCuiITcCEOjqsXfCr/A2Oo4Bm6KiObhBMlrAa45MPtM6j/Nt748
QNmBMOaGxaAW3pY3fZcCqAn53Ab3XBNSngLn5rLG9ks4pDrBukLiJiC5LGe/+b6yvKGLl2cB9SQv
mpvfmP6IEMiI8AnXSHy5CYp/3pfQEOVzGNd/jd2SBua3rWm1zpAYByT7xKovuXuhxk8Ebo+tMLIV
yQUXToCSC5FOtp4dALAxMWIO9C0y0UAxNX0N/PiF754uC9rVB8FWNCC2ysmLYmIezjhXMV86e0E+
TrX0n9/IALoeq0E/1SOT5IsuGPV8YJQuzItuRj2JqYX4xvdKSGweB1NSF6OJGFDDfbxatN5BZbdi
bRyoI9OBFBX23Z8ZzU32LpzoiWKdCUQXvVpkHq/1eVZZY8L4FxJhSYMQL6IwVhqX/QeS62ix2ItI
Ov8lzBweHHbhTULHwqoUi71dSSLlpsMxGyimV53ovwzTRANv5H6TIrps0Qcg+e4SIuIXUmkXoqEf
DTnMFHiETVeWqha9SnjO/IfnpATucIXyWa7WVBaI03YGWEnKItenZKMQBdITWqgTABkEhC1mWEoN
sVsfexKVaab+02YOqxyV7tm4vxe5mnNa3WzwPrKlcFBgI6ReVwuCv9WGYDJHkqcRWtdd2ptxbDuH
HPLwyhbwljvemtIuMyMV/ktfG4I2b9xldeMc4oDZr7b7xBv4pXYPt30x4PDTX4Aux4JLSwJo9EAB
dYTZuNj7e3LvGPiWh2lMZINDYk45ZcDDFTDzO3y39KXOAD56Ih7AfkoVcz5VKu/g0WFrqDOP0F0N
86CDw2ys1xeVNTe6wRVx4Bd2t//WPWWnzsJnXWaMt0txT57R9JptJo8C7EcMlPmqandAK3NvyUDa
kpk9gzNrE71NfsYGcwG2HCAUA5L7l4Raj+8GacwKSnSd5WH1YcSa6S51jt+XHufCn5j1s8RXMMRD
+DHhQVw8d8rvOxixbfa77Zw7vx7IlUl7+dyR6ADbLtwQtvHLyM5PoFvm44BLP1dEXNQc9M3j5lJQ
dHlMTnds18BUXwAGx1UA1karvuwUBbkEB+FoPOwEv8bhE6D7L05iTY7Ycx0pxRtn0Dyyfp9MOMyx
dxD/OkPDE4TuWt1VDXFHMuc/FpKa1+VjYASHy3ciW/BA7jPVebuACYUWxfRHNy9/1kD5oI98ms+S
gxbgSjDhiQTWx9Rh+7TpOFYMkRyx1BaF2ttfiQ5Z/KdbPgK/UL3MTUrQDbgScrSQCKfLBoTfKEw8
f28V0ExsAZo+HE+veI4SOnNm54qOVHfZDe27pBWzfTqRFFJCu+kfz5dHUy1iG0z+JyntNZSI7LQB
8R3pda7sT4UUnm+NubQUvRHUnrQ4kNZTeKtIIfgGbhhisFjeZ9zo/9hPnC5hVkHxWsfB9qMk4TPw
gdJpJjgN5pKTCf36XH3t2cnWrmpR6u/viRJj+yzZfMq0Y16ueJe4TN2l51ZhnTPzaRnqDbv9JdoP
vX0EdKHQ6Od/uPwbTVTvoNWknL4PlPZ5UYJa+UKSUUn05F/c2vk2bxBMqVryYSdqBpaLZG3R5VCj
iI0s0NqTuj/IXtJM5yTiaB0skJdMoKZ5Ww40+2LKYn9XLXvtezPesLWJZJMWDL2qMJPEhJhU0bYd
8lK9gTBi6OY+LugNUtHIqkTbL6y53SsEyTJKP+Yk/m7rkM8b79LE5qIkerbURN7p17N2D4LRFAnd
Hr3zhghvflN+7sbCb2dALxmG8qk0IwQbSJjf8ZF7+r0iMbNl+hJn9MYUOIjIfiGYriNzz6opUcFh
Ygkpt3OIuC3Ryilxh3i6pcsROpkKtKLBQ61Z+ooqk1P1dmWyvHeovmmIYL9fxcKDfC4U/gcmsXrh
BvNqS6mUc/SMtFR5r4y54KzyljJDCnTEK/0nkL5+aENDuMWYrvtIbqCPRgxS2HYqPatyhDTN61Ue
OTzvPONn0OW3aUyzbNaTJcFTrSv6kyHUPWDyHG6JgAwsU5vVroAKwqWXjHN0whzoN17Q31/0m+4F
/oRnIOdXE6MYUHsw/GMT9xQtWWGYPMIaoiksHI27w0PsgH6qDYMC1MoaEUea0oKg+y+MW00mPefI
TtT4iS5Kaa/uoJAqXNiXiXFPrt7WpbBkM58KRHKfgGfhB9gysWVNecn1IT2L1uN751OCt9XuEZ7+
bFXZWwOmb/kpbN7WIJwNmdIkz6ekxRI5AHPpEkVQbEyiPeXxGVw+ztXvvUdlJcQPThj5JtKsPquD
Xh2M4oCmrDmSrGz8LD2xgra9ZjwQWPNCjKYHpVX69Dz51dCOk51sZ2B7dgOisxO9p6r59j9cxhru
PHstSZBlSGmgJJWW6qcggPRBgRRxCTO3hk4UhXdML6hdR43rQrcsKkmLwclGrMV2jQybMQk9f9Cb
hmqBUVuyH578ydyIWOgShyjY3DgFBcQdiRufwiMgUCSEwbeYOq8X/I8lExbp+P8Y+Q5Z4gCcFIO/
7A/jDyq7EZRSK9s31iMyf/wq0YZ04hVgj2HQAphAEYvh9mmRSGPeaQA/j2lPwTaomX6FxzGYUkhd
6luMW8DH0rvmXORY6PWxnYF0xgriM9JfaysAK4ebfSL3CIQOgSAX39EixY1iASbAYF4N1ydGYVCf
IskOYILqJQg3NKzf8r0Em47WwB6ANuI83AOe5l6kG3ZrjCawKpkPEsIQp7dfL2EevLcItY4O7WzS
12+zo3A2EDwVx0Vr4oFSeWgZ0bPpt9Pp3QTw03KxRsgS1/xhn+MGmsaqPFrhfUNxtCAhE/6E874e
vYha6iSaQFcDXFl9Dtz3CywkvMdG9VmP+jPZ0JZfSiYM7m5T7rui6hW88ZdGJL7VU2B7GkNe/QnK
rs2AIYW7IW5c2aaF3orgTFfHbB52BwXnTZcT1yQZ2NTH1F/pS2Fyil1ZFzvJquMemiDrB9YY8hhN
gsn1Ljdi48c3BYwHSVl2prwJjIAcLEH2JUv0ajP+y4FVO8X5RqhXfW8qBqZ/nsbIAo5rYu1iPu7w
w1DPKHacnCAu9eBCdZdKFeGOBmTc6obfZdWgTxhK70bvrZv6IhA4+0PetkGjriS5TbYgOc05disf
/+X7Sip5Dyr1vD5n3OplFHX9BlV2ZOTuAUJ/mIz86eQG4Nq4NfyVuKg+WnfaPdJOzaZ9yU5J4JH1
oFWr2KfUKkV3/meaBONjK3B2095x5bLcXrWJMEsTsDUfRL1oJbdC+1fGoHDiaRZq/SE0iHolbyFG
Ix07nGxW11wIrSr+XbT+LI3w4Mz4MpTCyPxQnOqe6/I2dJnHF46uyilip++H72OF476gycbpFlnV
0JBTarh4hRYpr1t77q2n2yiBEOVI7buGbk09vcRkPUIgtZNBXsHrgLVmRyvF8EGB4vgSxTxunkmr
5ra4T1xbdcuinwbNFNxcDqBQLPaPaR3Ks7Yv2pzu74z58zNMjfr14ihPbTKt5Hz4o0oMJsrhFV91
s+a/PJFOSHLEUJDwzijoEwqklDPtT41di3c+VdKaRFvi8Kk8sm5j5WhmL5ehXxCat5yCdcZsQs/2
PFq2eTx5ESLlawSHg35y21z0cRNTiu32OZ9+p5BIBWngjKBUm5WojVeDF/qn/eJRXnGoZkWVmq3C
+COMz2GaNQj/1G7HsXxGlOlivOqxThZDqrz86K/Yq9PrihAxVlaSkXjGoECiQMb/MXKh5lhGFYCJ
mwtyGHKY8YctOOWT1Wg8fNeoEn8XvtdrZY9ov1zSvji/Emhnl6AQfk7WZ2lRyQU7KjtPSgTuAzwK
MgWl2z2xvqgLcyQo/NZPKHYrcINlk9bnBtYdKB5TPd2+hMWohoKTn4ee2S0I2wcA5Lr1r5vzuWro
JZk0bVizfYnqt48GyRxXcpQiK49un512k8eYli3sE2bCA4H6s2pmFAhRZ83npiJLxH1PfI5iZFtW
xgY0ebfzMcGbviom+4F7RaHc81GcGdCnMkhYD6la0YcGhzqPAbIIyG+QtN9xireuGUfe6Jx8UTke
kiFCewP7RGZ8ewmad1FIr4Mqkqfsc0nZOncFDQb5q3W+brRQxy8R7mutWLnVqVUdnMC4n+jtP77M
7FNpfAxyw4oLqyTkN2bi3Kb5kWM5OZYMWccVc1fPy1we2Itm+SjOqo55KS9Ft+jSurvnnsmhEYyS
UuefFmfTjfdUr1oxn++QSzXyhDRvEr0Od+BVkqWNsELyKJsWiTv5EAH6WWmQloF0Z4y5Kl5DCyzC
ycDuZQ+8YzFC1IqL4W/ThrnNG+W3B9rg6lU/XQ5HMGic6Dj3aMzbAX+f1lY5xEBji5qmm9L6kckZ
mjetcDgDK9hzsu5EMD248hFJ7gqCjFQjehsxDmWEX4c7J+Wn6QpZlA7DUx9hkCkvfH30oBrsrrqH
HCM6li81bDCaTkYESJ5UQjhNoJvYhaF14HbBr7+GqZkKTkwlR4/S0thdIruG5voRkdiFEE2T994I
HwKCuBIk+rgwd/AywMS+CtqOSr204Yd2ed+TdAevLO0pZkXJswjLLJv5z2A/eWNA4gulzkVgjCQW
WBxnc41ZKsOXiR9T/Q1lPFPz9+IU86rvS7lTwzLk65nX4sKztdd9wP5GCC8TXzkd4p7WeZGyBGpb
XXWyh1D63HbxripCcXraVi9ZT4zejz5nLc0T/TlPCkq6GV0M25CPiH3btNpPWR98L79ifJ+1zvS9
bQksIUllEgsEYpWqW+xFxa/zY76yGyAlRsGOi2nZEkLVIjeoLvqcXXYJo523Av9f236vLiNd7cXH
pQEdiklAYUR95juNZTuprlmQq4pErkNU+p49o2CmK5LR024QH6BpdZOQnI8yMS/DjKGWi/id/uxQ
wDkADlUC0CIIuiDiZ6Lh5rLAgJ8ksrm2KkgtqoDvumP8HQKIwybUePoo3liK8oZzZ3vtpuQmvi38
/XjETinrQkTE9C8hGyHuhIBZ5AYpwf2tDaEHmQxtgy/LfMxFT7DduWW/arMqJ3YPPDIg/1AyNK/S
tnq4rA3zyGnAQWX106IGQDyIH304yevgmAKLy8H8E6aEbf/bkY2HtCl15UHE1aPphzyus9rXSQle
kgCwh+dTKVKTJa1f/4AuWfNUebqEpGkKIOzbDDhnudSV5iwJSc2bHbv7J6yxgg4Zj1CW59WhHN3d
xqhuvRUdH1rqSo7tU1rOJWvcNAIcpYKAOvzbnQ9+A30EP2JPFrjPX23PnVXFACf1YsGltcCzQORS
2TYHBozligXsPF8alvHI5fKvySFnTMqA04hu/i3L0V4jUXIH7Vex9rQ9ALisplUoZimVpqR6L8ob
hKz15l5qyWrdeAyNcOmD6TyS843M40Z4Pn6ce6NVjyL0Ks7RzPwsv1r1FRb+V+Ae4z+Z/6D4gZDf
30xLre5i9Cdaz7x4Yj1HeuiftL8+w6qjSKqCF/GHvCa+n53AZjnxeHInIBSMJOOCNBDgiGG26bXi
uCvxV09uz7DSFj9aawuV5jVzfR7p0lTCrzrXPzbeE342YPDA7ancN7J5N5/O90Y2fmnYbvjlsQ5g
i0iRch9R8tyaldfNxUormb/LR5drSsDUCly3TP0toBA/MMZq4GhXYv8LoxAJ7nPkja/6dYI5uKoF
WCc+U548FKC95X5R/zvzGIju2d81MXcdbUp2kshj1pQoUf9M3Im+fSs/EfhppkgjX8fQPjP/r7ZT
22W2d2ScrM8tFtNFv1Pf71z511eE8Lfk8zta4EfmEmXeNepQt/EJbMbhHLHYTdi6IVHtQUUY7BtA
E4AbqWwsGoXwohXuJatkEr84jq0KM+I0CXvisQhni959Osz3gTV83JNmjFnTJSR5CcfCTdqga9Nl
gfczQbMgv2tDuoIkRHSLz8HeMz6jOvgq3q/RoceFVkSWKNDw88BmVGxP4bv5uNVOlOtrZtdBkC6i
08Y7JiYkoZvjy24Bw8DOPsPTmclP4Uz4yTG2PZR2IMdVR2B5XPv4dSWbc0Mf4cTFMpCLxihgUtPV
fvlt0swu4UmgNyFyapi37PqvJGYYt78zJgPCCtLcRcHO7XUlRnW6MHrT+HmGN1cgtWcV66wTESDW
5n3Cg9b17LwCj+8T3g82FCAp9Ojfwm+68rxoEAQH1hE1NHSbiLzuiZJGjVv7YbSFWLVgUCgq7Bq0
iqF9v8wY70qZwZJsjLe26BfPkQHULiWkC8w/V0qzmjP3OiZZqjyhtY2F9tdHq3v8oWl9M7/B+VaJ
5wtYSQV29zDFj7nj9TCmjxOOWk2PnDwjqLFROpx7xpZbrIGYWuLEuw4VhO9tyi6cMVgTSvdQ8HnY
kpFuhECN7u6WrNeeqKJ2xza8NFRfzNJxZeWZWJK6jxT8llWI6R096tcvklqWkKm3ANoaLx5kYaNp
PrdoV94BNNvQInQDClqxZNn8udtJVzeH3hVCVRsiOzJuSmd90BOB9nL+VxjIEaiuyWR05OcBAJQ1
BMO1ytUSYIdYbUW4Ir3zBPwotXJqAZzuNZpIKE0/uXCUNVFjhH7KULhpk5yPw990yse2Gg7V2m+V
NSp+3apiqtxpgvX8n3BmoKYEeM+CoODXQjd8rE8j9IR/htTl/E+Dn41sDPlhQjd/f4yRvyDt4LkV
2/9o/3FF7qZlg7UMeGW+0xc7A4tPo1nLFJij2hwSyKMFRRgzbYPSZIg6m3HkAImjhcFL9Ru4vjpk
mb9hqkalG1B5in3gs8gE6G6cqOpHZ6HvP0oqQ21nLbA7NMsmHCeIECh2+dcXwuBwAhcruhI8iH+I
a4W/qmBDeR7+b4wNBACDXBn7nxGlPyR1l8hqrBPFbOInrKOSZ61e73LExXMUYITAFIlYs9lXCBYr
pCw1u9dzuaWyj4YElLyF2quFIFLml/19aevMPX5FE3FSRk9j9TnjXz8QqLmdnDPNzs4fvtEj5o+u
rEh+qiJYhuoDSiSHq/KpxQ9tnSwtor8FWEoISA/ahW/wCxU/JlxZ0FP78pLT4Lnjqc/WjbBYLEbe
95JebzaSwQfQS0lRc+XXrdnuqa1HO8iwBfB0WqYwCtGJCBeBPVyVvCRgKoYl7d2uZVljEuLy2XqO
hRGlEewsDlmlKCbi5+WByCpUmUE46b0Iq2ByqTxXvAWTZGvnKwIQulqHZZ6fSxFc/LqmxteKyoyo
GVmSQvJ1ddwmJrCSODtuVLwvHLKO7rckmoaPIR/vlQTLKatAN+QlnJvROiibInzYJux/+bQiptAO
gOO24wEWM8e4p/7eYck7LVt57ZV18mCrYw+76bfB+KSUIrnhmYhbc86+QVfENU/4X+Mt0nh0pDmd
1P7ZVfKpdj4kgdWi7ca2mhoPH6QSSJuyQlDVEjRPxRqh6u4KX/d0GOdH0JJwobGMBHwKQWwVUFSV
GEK2javzqlsPsnmOnmS7CrCexAWV7s3ohJhM20lQ/hQxRkN/OtpRMJkWG19R3Fc84fnQngccslmi
vTQXCYVFP1FS8Z03x/YGDqwhJe8G9y4fFgSjXOaM4iPzZTp8bRh1c/Z+lNRYwgVHq6i+p4MdqwDl
u3jdSDwBtW5PfWQXaxGgDMvbXAnuSPx1iPrsfd+TAu5f6ynPGMMBKALxlURFyXsMFZEO0H0l19qy
g8n+zutG1KbCpKhLof4wLkW2cYbrCKFxjiNTf0Ik29jjKHlAI2WG087nKqDqe6j0/3Iouh/qIHTC
pm0lpnxc8liHi+LW5LEmcVPagYgnjVPv/QeDCnWiy3MhvWXmQC3oFNE3jtLShaFiGgoB/a976oSn
BaQjSPOwg63TQKChsPkG45o2+m5OkRGPX8WipV4iSAwXrg/ST8VNrBhRU+uNdFbRhcJrGue0chLV
31/WlD/6h8oD4EeOAF5KQKJKtFheMyszvWU/xEA8Wn/ez0ZQ7Yx8cjrA+DV4ekm7nxGktw/jC+lB
Il+W++EVD/E2djCJzo+fI09xZUlJPShKTyTOEjiBWe7DZshCGwMdrtSe0iX1wkfvyVLF8agHk1Vh
YE6chS7yLksiE0tkSWikbFOrRxdSK2t8anmahXtL1YKmmXePHUODxjMoDDJh9A0RSm5iJWpz3pas
/2lt6w7MrM/tiGlC8tUAS8/bKzpqPGjEg1Fl8r3Dh+gTgJ7+jBUUnBdss7uv3TqpKRdfoyhhqZW3
mTvCdvR3SH45J6umDjY4elKmfttJCM1rJUDZuJiO8nG7orDp8nyuBF6BHdwLT+ouGmUM7TWpn1wk
42rYpmaX2jCG/SY0x7td91/XstcjnzVYpjmcHN/wO4RUtJ55TSwfxBqQ7JZP80Fk+3UbktfN/s41
Dl08Ub58GkF0CUT+Bow8tPMwKKIiWm786OpLg0uUdFY6ZYvK8iAmZQMTeH2wf42cb+9nT+PmPtEt
izF6rBpTvGvXhIrwIzoiDIGbPr/NpLNaTITXOqeLKClZctR+deqqvGzzON5n1NZQ+f590+hr8NLf
cFESaFoGhvOAopt4Qg/BMlZ4i0TcgqvSGt9e3hG6YV+wj64Ya4YkB6X5lzd8HK7gqDHVuzvacV8i
bdLXyUK4cOxB9g8RZBS98FdAz+Y6cEtdLDOZYHttBJyb7bcu8meXtYvht2tKpPpkk/HUezL71Fn1
Hs0GzrTyY29TTs97D73/7FgKHxRhCxopGYfq0d+jLJy5ifj3db1ptzwL7fya5LflealaRvK/x/hv
ewnQBjaMzAn0O0Y7gEQVA4HeJK+z9V1PLOytwnc2UovNjjoOVHP/mermG1yERnPP+eXQDAKjD9JP
e2u3FsuxiykMxac6HboMpJcrWGKAeYsqungl5AWaFnr5/4GqcGOlJCcqwVO+pQk1VeqYnFAr8Nc1
zRZEemRmRlsHMkHFjaWlEXAJPNtl0RWhirpu2PD14XBWXjR5hnWCdSPbUO+nCe+mcN29h+8olezl
VnzXlzHfRSE+0H9Y4cpLHirLJmIp4pnhlZNMO8v1DUSlxlJqFU/9o7xKmFg4+ev+JUU+3N3Y/XeQ
cBhtw26d1+169JHvrVWaFNRcEwysl0k6yBpE3lFXDQRhokgMprt0fkkNNOXZ3U2DimyWRM1SlmNf
4BM/9L4eRCfZrWn8Nc2mVPn+HWAB2G/HAQknoGt9O+qywHuuJtv14hX4C0umqG/fE4TiqPZB1urK
OTf8yi8toFvoT62QY6TVM6TpVqM9e5iSLE22CVUh/BDMFmYXwdGdrJ+AnRgl9+jMB14Bx039gXSX
90qiWs9DzilXepDXLnV0hmdkJ40AaX6FNSzhepqVIZpN3e+zI6qENo5VJI5e0F7EZTCYXdsyoFBc
rSNZSMclQU2Dug3cVUGcf97/TgjG5BX7Ks1iFzYdjtIMIx5jE4mN/pyn1bR9tFjRwjHdaSNGHHws
5M2qcZzMTCtXl0VGChDZTu4cx9dTLia9wYXZdQ//9CKQrIcGyB6hzae4mnPUuPVpKky3V+V5BsgT
zhoKXWdRdoLDWSufPlXYPtuzxQF/TRX/R42pDRVITEyw3/mlb9Dri/z1pf3rc5eLcGDaz9/LrKPU
ezyMZ0MQa7nHBogy49bHNOLfe8FIOHVQ7hLxrUHPGOgjZ8JC+pY+C2QwKRMM8XsGM7F80DrXHmq+
0TM8ENB8K7C3SMOn7kCn4DqTBCYKJ1CqqiW3UnEws7G6QNHHsn2vDVGzavpC1NCT/bwDH3JJrS9l
bLw2kko4dadIe/TzPaUAxBkmKWPe7uFRLoJZfQoKu6Zo7LtE2LG2Fb8uYZNTaFEdzq3V2g7gZeM5
7kjDpYZhBrEEys8Xb25WaVwAE6oflKYfOIJVFo9w4DQvBJ/h4G3Z2GP8Ij31GAc9Ig3jcIfKpAMO
pobIisdqcIFMB6aQwaa7ndOURvwLnfS5yddY//A9q81i/ugM4uDFlhi08+oWWrU8JOpFjKyT9Hr9
uTUi+XYM5pqkrA0YZr6gW+JWKlQUr2SVxcSuMKSCyRUNrTRmlfsCg5nnddTGXvuH4AZWStwaaZdd
rITtPxF+105fbmpF+Z8xhsPQ2e/DJVyX0U5B59RvkfSl8aVIK7MW9gs/quURAr/KmvHKn8xdJXYX
gOmIXMbcFAzxIWKaed0eMxuyVWOadveSYEA2Ri95ImGCQFrvHtSxRvSce7qyos7d6upoVRlkpqMP
LRwNYsfgaheGDp0QK4VXNxEBtKKqmX17LefBZYNB42S5vweRUkpK797JG5axptNKKmzdUqaEn5QB
U1U04U1pkKCuzF7wu//47UBj4yrtxSk+ljqYdHWDGX2AdBuPursAI4jdD3MzbvjOLoRoAU6gEdkS
sL9LL8MlcIU9ZIMBJd4ytAbM7OizzaaY0TVqWnabNF9g/XIk5fCBVEdfh12uluskLvIPu9uORhwB
6W0pUCNyUuUdA7njZ9+nEM1Hme10lRroKVnSK9+ShEuezqOmMWO/33sOWLdneX19JEyegrfIttoO
nix3FrvJhSQ4CX/LaPZI/pMXd8qpy50XVneY6G4197R10tnsoaL8cYVVtamZ/Z2E84doahNBaeiW
QoE4MpfNZSLdkeVH6jVf1J7b2Vtn3x8giRuMC7H73cDb4bMDUrRflOR4V2gCSBQex4gLbH40z8me
i0dxiOfjbi27XsPwpGgeOHhix2F4Hk+uHF7ToLRceCuUkjbIyiHWzaS+SrRNneY+nKRVYCbDC63S
1JMeGEkT+BGluFf9RZkvE4nxJUbKGFUK4FUM4x4FlXtgDgIdnVakEkByRmuKRF89do51VSTZdi4l
BuzMlWBBoru9Lz5SeMsADtLK4FQbfyCqHB1NC32o6vQDzJ406vziUlVcf49zlg5ML9ET4qNO/Xmm
nHCBQ0Fkp6LrgpiJLqbzrVlP4SZ5btf/DySl8jrUJ0Weu5Tk4YAp5tH6Rz/IM9aWxhrczUj3YB9T
d19ap+wZLcrl2npOiqorW950OYsJB6vfjvXPt04pHqv3l4L0DM/T/xpIjQkBmxcIGRK7+T+p9cXL
RibM0zT6MZ4yzvIEemEa/oxY4GhM67TykQmucddAIPg29zyh28TYLx/kZ23OIgTyNcYS+oP4L+rW
6urjC+rEUGdWjUFO1319CM5rg6GG3+I4aO2SFoj6/AqZK21TaOpVQ7D18oUyqZiaJIvjCmx5ly2K
cAAZXjJhc1tRoVkg58NYgKa/Jr/tfSt3O/KJJJJIWrYWMb0cBDSKO+zUiJO6YaTPbcOZ86F8yTP0
Nf0eBrK/Nk+2sLjrgDu+6ArnHtwkz47ENGzIc2Mr13kyYWzKFD2pe5w1SjaGIUTo+kc5pz6pttGt
8/+YMj2o30pYrRXWlnL0ZiVn88tyvsvse661BA7Kxx0SOfKLQmFFJcVBXXmqUP6ZZ+YauxNO8X5G
cBP6czQMYRe2qWzxk6LvnOjObG3dr7b7wN/rDQRVafril38suCEB0Ky0F3fsA52XetEU7R36wgY2
pNSa0cw9Y2Z7kXnnFGJfSVeCdPix/jdFJgYrmFTK1tlpEfomOOaxIPv4F8l0ka9MWwcvGeLYAEdO
Cl6b/ZGSPeRklKwsSxa44QO0am5YeJf95xKREai3IFjtfKTnZkwHkoaZvbLGkG7N9acoVZ6QE38P
yTwE9gWebpDfkdTiGaYVX4cAsQZsTce2cMJhAf5ooycBheSQXt22rNMJfcuxLR30k6d22g1Ia7Le
xg7CMFEy2Rfst1oHoklqg9QYhb7Np3ZjoU4sW9mbHAkZttTzY/yJk+jpTDSJ4Z8wK66h5lmhuVtd
j4wX806jQv3RKt+spShh0kFjhXQGAuulq9sI52ISYejhTCFzpwN1kxFUei1tTtyJo4ml3ZIINmjG
AZCjJwI2sueTgYBzbXSw50MwQZgQGSJwXRsOuQdow0w2umcyjec+1oObOJd1LiJcDDY5QixTZXih
Uy2BFmYmAVgS66ij4bu1zS1W1OAoo9G9zOSYHACAQBeRaU5e6POrDAVBTBNBRrCSGy/jU3TDVTuq
hmIA9fXq2ceGYXw2oV4jBkQKdSj/paHGaB+ZayT+mbzHbK8GZNc9wkn2X0FTNNPN66sgIOgOm8lf
/OnjMhCtZ4djlb6o0cwSQUupcNU3JDCb++eSbczIZCUBkXoyIAyJ5oXH8paEoj9HGix9UEuYyR9o
h34e1jfkjrmrzEO5N0YhtGs0EYUyzjZN4ijT6adIs383WX38P/7+4sMVtsE2MX87NmDAiQ8KSoMB
UFpdjmxjET1lmLVJkiidzhIQGBK8YOeLUJDuXJLOBxFemzpYG9kL0JNsOZ5aReOlUEzDneI0bt0R
JoZUkIg6gjc6gwfiUeq9yso4mR7rHkQmzGBrCu2kLXlY85HnIqRJeARroG6MMNmywmRsFR0+MXyp
Xx5ku2UrV1IjeAMTWVuDFw9i/1Iad1Z6tT3tU7n9x4EEumJrZ2XPygcN/wj1S3AY434d9/muvQHe
675W0zsQJvADoyU3oKJG3l4qMx4Hv4q7boQ8yfS7R4gJ8Jw0B6a+m72f0Z4PpDPj5yl1VXxMScOd
Z1ffrI4HZ0WgZH0a2TSvgcXTuUFPSD7V00nIxVpcGD2RRdB/1i5wKmeEjPwzOiUccgJIu1MpTe7z
ZHLCb5UQfPodZM27uADx1v+IwN9HcUtDNTPxKT18iy/ERnP/8fdEg5wRzpaT7Vkczs9X9ujryx3l
w7TP9wNDdhpHw0dtMAuvkz557mXUXtoPh+WAq/CR5V7DBBdF31Bxid/shaIBGfW8jBrQHqjbrYFr
2gY/ZIM3vG8WamtDuhlBeD/yAO5P3M3ezeMRIMIUyK5O6r01tLz7G3Pl1vREnSycNTbCG5MvOuIe
/eEzEdvKbL0ZucKbrhKTvU75lo05CK6Qr7a64gQEM6C5w3iV6WTrp1L8tNwiIlags+E7ksBgMsPi
IOvWlOkFGss+rL5mSaeIKHwVKk50XWBdLUxNQGWHmSm69MZyk7MRAPNGU6eRd2gYwqxY7xwEzok5
J/67hWguULW9UCPI9cuAiNKQEvw4sMiG7yyiWq9ChgLufNC7tVojlZeSAUl5oq2aFQ8nCglF+6Gv
syiljHsUMszj4zgWY0Zz58NhtLnYX37wfhREuS0VbrY+LvlNinKiQTaLl8r7GEFdTxh6WBHMConx
aQy5z446/Ia/XW9DYPbM+iqSxFNJIpO53HRCOOktfsmgZd+hpvOPxasdSgEQ8aU9ZZD1/a3us04I
GUpr9nLfSidUBBNLyuRGHeqIm9WWZMWAT3TPPjZSQjSNP3+Xyx/rrGJmN8G0XsC4gm6GCrfYRYKG
mJfZSPZetI6/2wgKt6dThh/ij1E1b+SqUlBuaafluqhcMKurW7vjJW76wwXSEeYpBns9RSWBt1xC
BFdDKXEsts+SB27WKnVGEZBmfo+n4EA1WQU/D7zvES7lTeW/IeZ1WfdyzdZEgvoS1bKUCvbyzoy6
lt5knvnwCyAurV+2IqwlqmNxPWv3G3sXCRqWwIV0mw+AnHn6hmEsS0XY2fduxK0ypx9gZCi8jhsr
vWWuPoxTNIMil1tqgIf991gZzorim3Cg97Y05mdghDlXzp8SrAtg35YQX6hYaWSahiGPzz67/e+x
8P+mAKrs3iS7A37YXuTIK01Y3mtiwP+mDpGzei4BshJir11jTIu1UKFGc4jLd5IGuDugAjxkANzu
liWfrQbkeh3DtMvBL+PDqpyARLho6M1QO4PD/WSmnruEds5anP94Dmrp/Jd+HMX6bymf/C4EUI1t
ZRem9S5KOu/qXZKvamGySrahw++mkQ8W5kBeEA/T/2EUDe8LWxxa2/rwKK2gEdKdGti2bHLCCVZr
hMJsLiduH3TLDCPvWCHQTiAuG9eIOFm5uulTfa99H+brrTcP/9n+Ftxtk8e37AbI7XkvkmTkA7R3
GuhddS/FOI2eSnzF8kbrXKbEjnIPvvkQ+NL7RGRnqbrkC5kSG/m+tpWd2Wc3fwZczY4WQz05GJLY
bxjTKlKMwrhk7YQqUBNxUIuaVT4re5KRAQHNFmVTs0sjFvcsWYAh2tMdsGQInppGIzgZs69AQEYb
jXPpEQUlXVoasGKkkF+RfPbVOj5Jf+zOb4Ok+J3xOta8WSfDTCfOLICHx8RxOvL2jiM0YHOtNSbs
WpwV4gSs24zgWNkolEGNZyCYcfTHUD1HtjdF9h7HBlRWquEiLI6tfnFk3eIgcWnqFjeOn19rhc33
JvM4KfSxJlZ6Hvz8bLC3aiKtF+J/fW0ETF3GJYFiAkDwnlFbZH275fl97uHzE+Kpkz/Cyn4omU0B
kisvMBOs6QDbhm0QGpLmjGVaxtjMzAail9TB5sb+/19iL2H8PhsODt4+JQprVIBMa1cKyIFLwnA1
kwWxDjUC5QKcZYKvw8fnKIIjYzdHwyd89OHbNZfztCBqVFA1HxZCCZH7Kidu9FdIA7DmnhPvY0h0
/VJxUAb0rd2TR7oLEoG7s//VCBCNhIWfI9CZViq23piYpy+eDOj6zI0h1JCtx0qv6qPEHS0CTx+Z
+QEsirJVXoqr2PFvxpVmusok8Z0SQPB60tsnEfC44wcX0JA1KZeyFlRkl8e3ypHOWDiaz7lWN9h2
pyCjLMkqwYy4nwF4mEUvt/fKdLNVYDGzoec20fqXlB5vlKTqMQQQ6tLz/coZSofOIwDB30UKNB/Y
o4Ua6/QStI865Grg1ZSb87J3vR9PV4E3p9492EI37WboVSuF/tUVc+0KVZQXuuxIS9peblPUgh6Q
NRdULegec+yb/VYoWkm/uL+bkQmYYIJZYnXGkaogvAQxFo/aBVInCX1HyJwt/tyKBuuVy1ZDvuNY
CAFwkQ4A6Yp4JXJSIF4HU9wDVpkgiQ2rppQYAOU96pxQmFCDHZDXz6dga2I0aJJ2yOmkTvtsNhvq
C6dyhyHtuct5IDf6t578ydBnll7XQxEcm9fOaVTdDkaaMIBp/nohxkAtQ0vtdenkKhv5GQCk7riJ
9u81NPNkLvmn9RFQRO+1DrDjWrUPg6/f4wPSEGnvxZpTyrE00nmCVoKm/q+6VEjPQo1eX0t67U0J
isFaTvYJ4w/IhjnBFpgynLW+bzzcV9/zTZ0vVQe7YfLg+nDjSaHBzVEbev3rqezjH3arAzgqQ30Q
ZwvdbLWePlMWmQ+M/VxLfQ0ZPEiPV3K72If5u+z93ZrQs/G9che8yfftFVlY3dK7M8lUVW1kiy6u
D1CJrky2zFFxYMXrAQxewyifpojiusSrFMQZ3gShICyoS+NytwgX9AruoJA48Wm/oBF/KwiLTiUF
ayzSnlb/CrD4x6xg4hYb8qZ2sF+CrLN3mWJeDJGmGMPyFJQmeI0/pm7/lKokzjNFbGNdbBiYGmVM
H1aKGHzLGqqtcJxcAR8x+twt1W2dDPLkwYp+TNK94dhtnvMQ6dvikbv4RdwX00eZKcTj9Y4ID5Du
gyJV9MJMqK0S6v4dlw9ZocDc0eYBpGY9aboDVomln7LOShSw+VEQXhDqFPYYg1PorbBl1COVCBGj
R6fcaIovftCMwwtsVUNNXYHOhMeF+UGQVVJ+ajWNUlLCj04VYkfHD2hOT2dfe3C3AImbyvo6YEiG
4yNyPEzmUL9Kgkab4lZ+cDzLuXauwQaT5cbY4/4OVm0cDPriNb8GipW7qnId/JsAzqTx6mxHjt/a
Ok1k75Syp/qsvOUcUQKIUt1aZpm8EaftaRGGCpDcLfmAc8u5IIxbkWILHiZdhEXsvwmmyWcPw+um
fmXwUQeRieoDPKXMJWcd5tjUjSwdXfGoix59jfXhKMjpI2H1C7QfoAx4ETVITW+lfWYzZ2XdIk6v
5LZYx1PQHQE3SG8rTCragdOCKCVumjxzJuYT9isVoz1XEN/KRYaykymMTVQrRX6gzHcxCc5GbbDb
DraYzSVK2nxNGhZmxEMGufIE4TJAKWpPURO7gjwNNi4GFc6RhtTo4NdSNWMQ/cHeBkhe4YGrXJNw
HGxXMgCeFNYad5KOYiXhihzYsL3WOCraUSQrGaJhX7SDiIkZjXZUSJ1PX5aIUEq1JxVruaHQsshB
2/wVnobhM+wKsCZu29PEG3MZ5qiv8eoPhspgYsMHZEebym8xmfY6V3iTQ6HkXx0FQJIcweuyKhRB
PXObutzMsjRxvYohAaAjiBwqtuGP9lSv3kVvEwlFVeNkB78HEgBTa/Z/vFuUEalTeGmXZDHkVeGh
yOVZe35LkmsmiCYXl6BI7d312UuCxQcVYC0mRTiIjkQEkMHmrWGAle+ql/7IYHbE+DRNd9noKfiL
JrFxOEGr/Ipj65ccEfiGxndODnajyX7Nx1Qjs9TTwEgRV7zL1gfp4A5uc/ONpvJ2Uyv0TS/KRDP2
RnDRrM4x6xULWoUs77i7y2CfmDmNWWQodFb4DrUMUboXo8xoJu0LdPpp2l+Hxa+rIZALvFTgQ6RA
7CI6UScUy4wqvljXC+9c1Nj2RzPnUgq+k6ydZSLWZPC15rmvVgVwj5hohQCmvvMhkFcYPncGN/P2
7BI3VFGWhDFZUY3qyjDOR6mlFCUCoHHdoCCSALtmICSff8ft5HHejNcfTwooNo9lo8JL8YTkV0Ez
w69QYy6c0b1GakjTaUFPXd38/M8/GrjgUnekgOZXJcFLhzawGq8qjaVzaZ+UYeJpJ1LDvmTlzNTz
TH71cp3baTi2PSRgpGvumpVZk3aXTaWuGrn9JbNGf9CxVr83YZmfibQe01DIIwHWs2+dN9S5KMT0
tcCNe6xXOrMY8M6vho4SSDa42YeeEqoYBWNcmPDn1NQEx/S3a3AuEtCxP7XtfeSdxCdljk803Tvp
zHnnACba0Hzkl0VyzmuCKMyEtQLzv+ZNAxGthrbHEEz19F3tm6qgTHfZRnjKzCdZHTAOEXQWzWXz
SzI+7u26Bil7LMEmTr8pRxNo9IRMXNl+v0gCxTVgIimXA6Vh2+4/Uo0TM0rT+mz9bGcGXt7IEAnY
T+86h4udX2nOOxy8lwebpgqF+7mIJ775gCZbTDh1d4saGwT284fS6tjvWXT/xG4z7R74pgOpvnSs
DZeZPkK11XY8Sj5gdFd9BJZ+rLunWOOgprXaJu3FlfAcsYVZPQgnoM/t4Y9JZNWYh/zdXeUw72Yl
ac7yTOYofwAXP+DqwHkmVE0mEqt7flMRWLW3phEhGkr8j814id3hJcWqDpIsUJ9TKTrH3i9r1wNU
mYLQosNrLIPzpTIZst6Fif1p/Q3XEvEYrol/efAO/BVjbbWCU7OvdgYIR/RtcCMzgeaPQcwNPbVN
3ef9l1ADLCsyuAYOE8atF0qcbXYV4ya8ei2N7+JjX2ZyiCSMFj68JVb/AACnRCNABrqwkqFf1oiY
U0jnpigkd67v0Imamgz6lBqt1+dDadpNKMPZT8jUn5/CvSIgjydwMKT9IVWIH6GecTzaJsTnFt8n
us7w0BR3rIiPC0SaclQw1T9ezUVCs5OGjvKdjJi7HSXYDbmpQBSjqOHXCtM4/IYtK1RMbyQsQHkb
SkIsHj1T96lKjd0iPrfj9wvRCPElpCiX5fwIXBUc1KneD21IJYlJbOwso+UECOPTNZcNFEupLWxE
8T0qG5UBk8lDNowWFuA83bxCpacVsH/4q4K5S/mvp/InwrLEp0x7IfvAnHeLi1/f6bMRae1pvi/H
2Qt8UK5pXwdIoyk86aZTdgqXilLzwxsZjL6EbCRp8cbyKRFvkvmc6oglcRYeI7wc6Qlj4eh7j3c9
9zJDlY5rftBd7YayJiYVWekIYxhyNrBIDBErWQNi8WOOBhToFm5UVfecLazJ3i7etuw/GWqiIaXv
DleBsFCDx7780RR4WNbEP7jMxv8dWoCDqB4P4MHvKsWE1ddAqoTbzVWbNxJrGcjzs6wd07x3IyoV
h4itFByFZ/RpauvOGtpqAfBHM2K9VSGapUznfEkUgx32FMwBk/rGN+Go4JJTDVi7BXsV89FxTkrC
kHqggw0qwqw/XVx9z7t/NDDwB0qe3cin2wEazUqxVwPi/GhqwW5l2G+/6gDJJZyxlOCTECfkOQBn
94sbJnC5m5s5hk5FlEeFFA0ls8lmk5I12qIosFTuzWcS/u35vb04RCK/m5bahjGJ/tBgY2E3T+Qi
W1BTUD7otJdV8mmXG6XV8UMYAIO3yGFUm6L0zruAMRjRVBY6Yp3VgjA2U95/5FaEXNAXthdt1lLG
DQ8L043V5wmx/Odqd2nOc7XGEkWaWO2dOAi7p0szL9X4Nu66Y8/4gH5W8ZsoRnCY78ALIjgU5jTH
Knp3yIDxUpX73JSE7rQiyWdOaUNRHdRoA2pa2kK/ETBoHwzZWirDQsJNld/dSVTYej7S64/QWUcd
SvS0GTIB5JKNnCliB6d2zQhB8eUH9ljCHIqiu7oodC1Cbqz9nfqITgAwKxVpqOA28X+/72uEfeQm
8VbJwAN+B/jCG47eehaPDhlyGlNxPIK+iK9ow4w8sEz0pXRqG8mXlHZT6ldYL7btqVQlRL7t35Z5
vKcIRt55W+5ajrjOOpEQqTehBgPEnq8TD6Mq2f8nLAzXZgmrHmV+4MZUHTRuSGxBQp6BXppaDmpc
DHBG7wr6OFk10WvB46ON1JCTqUfkrjJy6IEamIyuNVd43RgvUZnTbqrBGQQJejHZCoINSBZyeOZE
AQHzqqnNkWyBz3jRbeHygCpoLW4gHde+pEfnTUWr14nq0HbwKvvzZ3jmcj6T2piOJt3utuLu+v0p
rBZdm8s6X/hRrtBS++k+5dlnYARjNWnzJZpv3ROzZhJz21N6bqlMpxPh3is+GKe7m7SzbZzRXR+H
3MvXsp1vNqcR8txDHfqyy4vrKIsloS68QbFEOpeCeUyOVsbMq0sr0iBSPDFwVUsQQ0IxUcoFANNJ
D5ocnFpcIBFlrFMXohgTR58+JrQ1I41wEBDMHD1WFUjvx/hb7bJxIqfT+JfdE8V9lrHP0RSTQL0Q
I+lAKtPaCkhrnsKL9zmt4Gk0/Oetd3vCSg+u773FVNhgHOK/uJvF9YdR4BGPuQ38jtQ5bObz+C4H
pM7csGL9xMQ916q7jsJFod5XbrhtaaRiBaxwETdvVtlxNDOCTj/uV+pOteO2ma/mar/GnUbR7YPP
1bLVJNvu4M2WU9I2FQCb8LGATAaxXTN/b/ushlad2WYMNQqEfB39OvMnRJ38qQmISlAO17gjElWT
iDxlXEfWKGmTebopqPMhySuUanpnvQytfhEqrgqsejEYIw22bjPINAe2+T7h4OQZXshHQULQVzRC
6UyZD7tp0X3VEg9piZ4juOCqSVJQ+Fx6bHf3L/BlOXpb3Yi9c2GADKADZpvzUG3My9Shntmhs23k
LOvDDr722GznChbVXabT5eQuio1loS2qnPdTX6eToUfD6Xiupl1HosIPGP+Pmb8u2CpFIpIkFFeX
trY6iY0qm3xte9u1r5wVC7eoYOrMAqk9hC/Ll4MH80lHpwDj5sWBeVj7RZ8QI4WKCRL+VrBJFk2M
w9iU61c/qE585/cBXRhx/LE2VKxP1+xxz07BzP8PZ8TxMAygYndjWOELKXNFFNFiIA+ekHfNLxID
Q7eeUWBIS+B0wrDuz+5VH9iqghYYOggHEfgNzRkIAO/6rsvezWYpgzuOPryYjDaNDZ1qhg9shSZ2
uPYQnKMqBOz/Boc7Cx/EDGSW6M7vvkHUx4z6nm8Fal/ntk2WmotynLI6X2t/vj6DW0RnGoPE7P0U
zkCGZjX+taL7eVQfcutmIcTa3PgWkT1eSRm0gPwcNafq+3sRaKLz2KrMNKJzsqgHJOzvaYtF5TgM
0/HKbkIc/0eD7IxlME+Wuc6LmJxwYNfPSRigcq6FOrC8X+qUS+3eKEwekQKl+BdekRFetOvP320W
Ufx5tHECk/32m45Si/cquiOqH66AKRk9o4R4PnGPC41wN4g8f8Y/FAR17MQY8MYE48YJvEXdGZnj
uDT5dXx5xtVTigxHzFg2fOMmf5cevotVl9Bc2TNHR3F3sMh2U4ZK8ATusdxVjhFXQK29EYUsFXpn
FiGPrqhGd9aqR9OS8W5t1Cj15hy0WNQls8D7OU0wRkzXQQDJAXvTk+hAgYGBD/JPphLvujzL6DQX
4SxFANcViUQNtgXXGMxvGZ9EyC3KT55f5crQuILD9MERNCK4xo6a2v6xxH6M5Wb185Fmkvqz2UDL
hisFMdKjSFi4hzDIUKJso9q/gd7SNPlNr6E5ffH03txZtU7VPlmEKmIpP6baM0vDks45dAi6h5VD
+WqPuc3ALseilycYpaEYsTTmFJ1DmcndUm9zslmGrYpDTqw6MQIJtQKlPNb9MZv2KEHs+xRf4KMf
wDFw85hgVMFUockilrSnsTFnQWew0i4/fYpjefJqPznaIgm36z2OkNJvPpnrslZ36j9dx2vPUXos
SIVbamWulliYuRvLv9QXoWsAU7X4da2+IlOxzmNo4yv7VbMOgUD6AydLsfgTx8hsnY8RUnEq/JAI
3MvZPMuxMU3uWLwK8sTTRouqY20EpqpfmzYBznyXEgJ0+/ov5hTr2942SwR5HRxcXH/DSyJjV5E+
hiPxdlh+C59kX+Qz/bVXFMICCqQkWUMeFZW+QO0MtrGda1jrBax0/wtsOMX+OtcvhvkK+1YTBKm8
UEeqVS6vvhgikcsU8fqcxItfMHgxgKU9Hiy2YOgT3n3lPdd2lo74SmkntxHFdQ7IjVg16qkiG9cI
RRgPyrSAQuoqFucXH2HQbJz80NLdJhSXREs4+oIVc2zOUrky3+lxBLOBwfxMM9J4dRv8sCgE8oYp
0ztnfaHi+TGXj3Nd51gHL58rZkt5HBt7GpKbEM9CPb+GC7Ex8dEIbgvFAeend6HOAvO+yKc+O31D
295RyFD0ffbspEOx+Y9OVej9tuXJU/ef6CVGWhPyv60MPdacptfJDJCFY2WNGEe41IT9bu1koYTZ
aBmVfhs8BqBwc5ewmhc3Ou9ZfWfucWl1Mt5HxeO1zmYGtVZQK1RtqAFbKBnLlO0CxNscEEzULluN
y+pscdccvhRntNgFpAPfdSVTLAXhbZmzffKswbO926JZomIsgmf8S9I3nhKgJDp2PjIsySApr1Zs
54k9f1xd1J0Hom8uIZgx4lKHRzG77/gU96aa0LfJl/1ty2+MiRdeC0lhNbhdcKdRlwO4G+1wXF6q
FB98bjAyW4L87LdNUeCSsJJymd1rVkyYMTo3zvCoaZqOwmqYQoZPXnlQoQuNXvveRNfgjsyZGKU1
bn0jzG2XliPUgqXiB9Vr9ibFqf+oOe/UwJZneJylavr8Q6fVIjLlphEjZ3aHwlHZNBrcQvKT/PJs
kOPEQjIuLMHOHmDX04Qmk4alON9kvjUmWKGbJDeIkN6toVhRqUW79CY7mx2V/TDpDM+otACKjIRL
iRHIC3Q3vyGQDjI45uYL43H54G7gn3rALO7zk6WvtPnIGdlMvKMvDqT1d1qCs2R1QhyZ54bSUiJV
tSkhF0oOLu0Ekvywqz8CfY/ZwtyMlW53fZoyqAOxlTbq6tX8HjtEGjTVy0kK/5LR3xAF+GLIqmrc
p/184i6MDhsQgDrNmWUTGWHBKEA3OOkp0ZZB3DbEY63BI6gmaaFIzjAPjzsxB1uZNcewTYTGcHWX
k+vwnwOvgNwWDLzOZyzrBcful7P4CAUGBgCrL70kpZFa8+9moQk71qpuOpuSo8QuBwM5+NrcM303
BhMifiD5ysUUggucDyEuGGx/ov18M8cn49Oi/MWG5XAF/NsiK2/fhrCoERh0CN5crMFM6QdQsQx+
SXUthcR2nDIaueKhNMvddrqd8X0In2hJP5wkAICS5LlwvVzvwpJ9YxtBwPRGhEU0sn/M0V3Qi6ez
S4lx+U11IBzfKm1Xcu+rwxmtM6/oNilq4IEwjsko6+NbtrU2E/ryY8bwFWMG1Cj/0flyX3ok6QN5
K9K4gN4afRW1nvt23UzJfIKzyJ2WCs7LkVAFKpjFOffU+5iYjY9ouikH2dc75fuvM77pPIM1RjBk
Bl+uk8u+HB3M2wETum0pw8WHZWJ7FHsq5Ps3Qn4IlNDrcFW01E60KJj3mZd5b/j/o08lItMYxjvi
iWd7/T9lAYNCMrYdF16NyOWxzaD4Dl6sIPCQZKv09vdfhH+uKh1aUpe8UStFwHA4ATcW0klkom8O
MzBTp+twdLcDhodimFzrZK8DkADoZXM0+yz94FDxonVXddjeAXJKDRCRXk5+f43nGjPbfr1P1UKn
HalWtssbr58nC0XGo25r9GJ2led/8bIvExNrFlFlGXNwi7ocJxik94OSIyYvU8JT09tnn34zOs9y
s1b0NeD8f/7RUVNm8FS/e/lV/L7Ia+U2A0BxeQxGjIh4iBjkBXJT+MHnq+3COFw94Hm8zEippnzh
jB8ViDSVTlU19KI7gvDvruaheIXjqKmysqvauJ7KnnF3q+Nh4LzfN/q8wKlegOlBuol6BT+/nd+T
yV+Xbg4JxO4TppXVLATn8730h4GLCpvlAUlb7aSRmRarra9medjYwyKpivsXqwO4r64oQqh72jV9
c7Duw3o54W1767c9O+Bl76IboA1cJ1AAqZ2VF3LOQqDynW9fESysDiwk6kkXmXTekDE3uPs6nWPS
cr5KuNi3ch74jCzFyFD6D6X0YlYKyVzMeMa1hFWNrMT2lgCZ3m/FyANua6clt/lyrls8fvUh+qMi
gBjmI6eAGS/SNmMsyQTWaJHpt6EHC6Bu7KY8rg1JHZJdpGT9uWYU554xgdL0O+er4/lmlvjRan2r
bs/1yx0cDzQkWueTPFq9Eudbctp3SXwMQQKYoDD1ijEmrI1HzZH44B6oEfWj4ZQhtDZnT4vUag83
oMWqoGbs4zoJ4ffysL05F1M5Oawd/exZ8ej/Qj/vg+6jcFcMLYVi3N2KspOXSZ7i3p6o5Dvt+vwe
lj73DOpdI5ffDk5LKAhwKPgiLkpmNGjOAdJ3tDNaXq1GUhvA3pS+QT9Z7tex2B+MsHQdVkz7OvjR
C3QLPcJyiSwf6/8hpovEjgU9ufrEFiFcH8PvG6fqSRwxtwOri+vo+6Fm+0Wk1h3BNA6jp+sckDRB
cTxEgyMtO3vjIcY70u9vAQnFKzpQT2Ny2gHALZlhNgx0ekLLoPfMyjQ9ZaJUEO7bw8K5bDhsfwa3
i+tsMFjsFXfIIEuxFocWFKsCMpdm9H16V/+7FhVPwpRM+qqI/Vh+zW1c2EgNcDaM1e+blYCGWGHB
BKyOo7ZotWwqLMNN7yPvS41XE0OHbHL/k5Qfkj+/lRIpry1Bwrq1YMAh09HFbiJ18mc/kvhzwSwn
0LJJnJJaQYSGC5g/NETogwMZv2qetjpD4ELKFvAarvUUNADGp45FiMD0kq/VqoCADpQJ9hmXwFgT
5WySf74zP9RiG+k/EC4WLtOBILKS9DAjP8YagJiUnG7uBygT0sfmAhCyspH2VszsiwxV4faAa3uA
fIYvpKqHb96JD8Iyjlx5NdUacuK4IP3SPn48kstZdaULGhcBPijzuaqHmqtajP00gMyNZPZse4Ef
YdhVihwvJYbRIp/pHnN7KiYhGGihLL8KNkMvhPy8kziNErbKL7uEjpddZbwHSOL9zYHWXWgWLGAn
ZMcsFgJs6FZuelRVyM1tGUDqDo68OK3HnEU2Pa3dmKgux+XpEtUubfeM2FPvm6ZMJegWyI0PvNw+
uUf2fQ/IJJU7Xhi8E2TcY191bPNm/J+pvRbaWUSsZCkH0h9tj+SgMReaH4b11xJ9iMQyJlRl7jCu
Ve35cQ2ZIHLhVk52ZQzzRNQ7f4MC2fugPLenrolG25qbpPV/HoV/4tmKN94ZxjpGrwmuAY3dROit
6Phk0Cigjjnc7nwFcqGZes9TLYWhsOxA6pUchhMB8yeGqWw3GFKECDVWHM5ckxCr0lpnXyWUXPi0
tlmreIzbXiM9gtmkjubAg6nTdrMcOZVDoat7DoIeejdWw7U6TdLGW764p/hXmOun3nGaN0H4w2CB
YVhdA0sfyjwVlMrKMi6/9rgvj6ZQAZ3Q93WY8C7EBDTy7M53W2ylpVyfwYIPI+aGknHv4Riiv8Gq
GWTgK2op5kgfsWzwOTKymi6fQhtqOopW30XraoyIg/a6pJBed8oONzL9ZLcS0Ul81Bx5amDwFtpv
YkfNB7CILIP3nT1To42Wjcd+MZ3X0OVnHJ7POuJ7qGhCyKzr/xUmCtlG231f3quHozntZd9yWWsN
0jO3w1vA5GiGyCNXQxD3GgNC4GOzzraX4vq8gUGwqVw/C5+3I9Lg8q1FyzVKK+pD+MDWXO7x1WLp
WRlu9/w+E85VgQMLLKOwkDzxZYotsoLGGGEDshZ4Cx2diXjn1rXIbygSJ5s+/qbDQeUl0B5IM1Ji
wUpNsAq1MW8qrEOdzXt1jdNEUQxkgCPjsABViJpRlUQT7Ol//aGi1z6qT25bH1wPfxhvmVKfrGLq
jGcY0bJteBykBQg5X3t7UGzzfnkagkefpRije3jbP6ditixcqpK7r2adGIsaHs1NYOP1tQuJZH0N
6xcnZs0alYqWB3cCu6WfYrNpFSAYCxT4Pva2hIocfbXSzSCfjGqemQro7T0s8MORUardXkuOvbXL
p03dLx2aB7oAYUg+TQcSRZ7uQKDCW3Pqwtlcd3bqZHac09kbSVjtHQqxMIpadIkRny9POd+lqVcc
1h8InIezOp092rxmxUZbRptmhJspv1Lph53b1LH4iDaBy1ESIDChVuBSfpmH10Uj30CWvmvV265d
sA5ksS/VyCEPEESU+J4cO63VvUBAsR6cFWITJ8qMvGAOPnVesy/fGZlvvteW1vWodd9qC/SGPXoe
kioCTGJqu+zf5llsUxzH2xVNCdFK63j2djFef/TvIeyTr81lKySCRb3zSZFGKeIT6bb0L4lu8cLD
SWn0u/BOSGGX3Q9MwvnQMX5KsKAHj7ub0LwZSyDv7SaUimzlK6pMFY4NCgoVw7e3qBhcvxmVeS1u
Of1yIFRdRyNyDP7wGKABtbKYPxgRa4tQ/aIuYTRuZDvVClgK/sEPkFwkF/FIkPgiaNRYh/IyspAo
JmMM1wTnGc0RfzmGVlJavia5bl+vodtIPBj1vThYC0eq70brkxfGhY4lwA8YpTpT5Pk7ORF3gy8b
rYtuDSyg1sZfxUdEm0Zf/y9PWP1+oHISQiee1yWWGSmh5HKM/tWZlJrGCK4/UpguKfRkU95QF3vd
0qN/xEZ5fCXNhrQ6IdtZKCVnaYmSZUOSfkQPbgb+CKjPbHTpVTGzww+v/W1Q95u5+1XGujVOPbfs
7bPFkKB+A8CbOIMVJ+2ihgSA89OID8uCqADU/7rpTkwwdDNz59WVlKLT2V+fLfLa7jJxRLi3Yzyb
ag04hteAYarpIw5onTsIRDzu1rvh6s+3vMglBy5h/clLE88arNpfw6XgrJxbz7/TWs5td1uT7OG0
OXqWjlM3vL8ZRnSWbF7sdLCFvZ53lDE8o2Mf5nlxsCRZh675rAfZc0rUFkHawI9O/8xrZ6t/EKE/
RM+lX4sjWhk8b96xBC/R+fYt3vGsFbwgk14/s543lMYUDJSCDSb53Ixs0TrAy18lEIG3xtvAGona
lQVrv2eKU9Gex0hVdo7YSoD3rdjT6UykBk5uiu0Ui0UEROJZgLWuselelnGWWDi1tXgKsGM4vO4S
2Q5QIoWRlzBu4t7U4cgfedom2DO9pP/8HaU+cTDnku1hlJfI1PR3fMiYL/GDb7c8Csr52Bh+775B
Ob25stEBROHyEPFw5hWh6ZUYMnTryzehXnn6ImPYJJMqILsJEYdLsphw1ycJGpOKT6Bdngg4nfCv
4TxmLezfi9csTyJ4VTEUVSc0w58iAWNQ1p4pV1GyEOYdl8phDVShfPaKt2zvceeRAWmi/28N5IGx
yp3FazrVKP862/VemQpdBZPKAFIRDbHFFYuTn5KjhkgflzE3/qS0/BYbjOEJmuAt+lpXkXf9pPzi
6aU2i8DPotvl0MeFEFmh1sccqs3B6+biEbFTf8vHB23NoCjfqohuMGJgEW0c8fbKu6ClcdP/L8m4
OJDaNQB+/tnDoSt5fFNoZiS48C2A1b85uC2AFT/g9fQpl/M82txIYekK4yTJm0U/Qf80NbzmQaUp
clvdzuWzZw2gb0JhzXilbG1uoPYZsBmu6UlCzrWlqJjNWS9A1UjmBEbWDAXi2MPi18n7EXYIkmPW
zLdwh1kHgCjGYHjFSwWj+sRIBwQn92eKlAQYg+KPCaQo4GDsJdsnmzxBFKBAapXpW4/1Z6ZQSjRQ
s4YAyT1lWUWOlsaKfB1COSlvn4rowxhnaPDp3Tk5OkwI5c15MpiyPma4CWCZm8j4WLKDWDlIx0T/
YmYXzHx6qMkyUYptfztc0rKm7IIhARiaJcCjbtFgYIdBjxKl/DL+KPvsN3OsIp+EZi8Ph4Uz/ps2
nlr8hDxS5BiinWM4sf7E5JVx7o0rcpWB+xZ9lTRL3EGD5MOmWQECWey5THdpxV5RcK0x0SHv0sF3
hkKYW8A9c0Z/+X1WXWeahXDt1IyodRzbnwe6kqclLnGUP1BVHOKT8Pc5jzDTOK//OSIa4Ec6Zqlj
KBTj88U7lD5pl1SjDe7na57iFngFzWqWLoIMMcjcZWQojvL/10gLZ5sDZ8XDLvZ9Ad3OfGWNHYo0
NsG8VvYwsPSPr4u7S65NrzizCqLrBH7/mcV2c7vjxCrYynNg6cye3iaw2cF26E/2vayKsil71DRG
2pr28+4hHfXIdF4ulcVrGyvvbGG/LEgE1vnw5kAQNh0FAaO2BIf2VGk3eY0X1y4/lncxSCGiCmoz
kA3CtcokuDN+jqLqXXFOq37z2BrNUfUShJYn+RFxFYGql2fIdmZRYvcGmKynj7L/gdlh2hQlaBCH
eJ7j5s3HbZua/mCbbfqFQXO1m5X/v14x07HVlArQVZyb1U/DWV4Qmg2iDQWD4B+VUZLeO6QwQ7Is
bR1lLVallPSGrcLFg65Vq4ga66A/NL06uG4HHviE5l6Ww4g+5nfvBuacHuJpB2DGjYALRMkPV/Nl
d93RXu0s9E7Ax1s1BKRrwPXmpyj7VP7zkWvezDfQ99R3MkPAwxi9+2w6Qt0r2yJ8e1q/8emF0Z6g
t94JV0DT6wJ+Nepw07xtijEwdSGTMF/Vr4gMZJzU9hyiTo7b3RYemi0CxeJ+nivTbVaam++FreC0
5bl07JKgPIfYICv7v9jS9HhqZ9DFFHyE5jqHatNXWVJufD5pNtIEZMhwq3LleK83AgSO92jgMmtJ
1w15YSbFi/AzX8ADrsOxuyln6ZGFdWqgKqIHxLaiVfyD8f+djlTVmHsXR24Glo1EXlG4OOl+p7WE
lLBIf8Qn9afIxRQtsliNQXtrX5ruGGzKTcZTl/CF7GvfiL5ANftcR4NqBQ/CLfCBI2H+MdqLFPab
CjrHriqAXkpU14Tysg4y1eyIbO9Os9fiz7vzG2ZAtr1vqM8O11DyKt6VwwwEEy0Lhft21I1FxCV7
INLydbYOQ+iO39Ercg1VktzimroxQ3SMG6P6uquBmKJT3HuGCHztupr7mK+Ox3GluCySDcGzIKpJ
KeGDZVzbiyaf3170WqwEtA0aVyBFkzY3l5F4+3rq41dsdd0PMkv3pku3BiUD2ubh84VIeStZT6A2
Uhob4K9Wt8bOlTH/BlbyPqjRWbbogHhxoW+Bj6HLFhvFvkmDgZ9JlnK7jouAnUKb7mNYnSh+Xl5a
qZRAXie213KOxecOXvEOw58PfUcabrVoNbhmwOh+bSEdjVtWMekSGmYnAspq5JyVjOOKExzCijwQ
XOW/oI41B9+fNJFCsGwSRHcxNJEoB22Cn0TmPEgEowP4D8UOW4I28+oLXkrSVB0ZPUhi/uSa6dQN
TPTJii568lND4e9i+aRLFzDbiOzxSw8BJGrm3VR+HNigDB73Butae3X86QqzdC96vz9hxFflcCw8
VxCVrjjstfkY5KHELA7LyoGkKBdp8+Nbu2fBhSoiSaX6fboaXtuGkovpxuv6s/2REMtQwGs96w8C
TgMCVaJPVi/gmUtFvqVhlFtGJD86mVtcqLiD3ykYdeuOEdYN20V8MpihTItUr0MTETppIkLzhvYD
/sSJzYD5hqo2q1sDpecN6NHcNlk86Zv9CHweo6SYpMEDPX5M43CIjbHsEz/6veUEiLsRrXDvqnVE
0XPfurOHJ6Fohi8/gJYoJHBpHjCZbKsvkayzgjTxrxiytBLWBk2cFkgqTXylKP41vyRny11nQJAF
ga3tl0nRtFFxKx/j0IkvgqS/wXFmgscAUZdl9sEQGBjltlFgjKzPg3MhNDmXZfRGGib9y1Jv1iHS
IXFeSFWEIwRNchczKaEfxawbRwHcrRmoaZL9MJCoZzahybinq0KtF/RQwa/Z17/Y8UERGySAdoiy
yenXqYL4a/2RB24qzzIYndZldYe4ll+8W7OoqqgHwn22ANPxRdl737tZJLO7RuMzENXGVXy605fH
0jGMgFfgNVnxLVe2lyhUIGoKSjHvih/sZPC9/qf0k70tBOxVrv83r5PGNb/NLTqeJvQ721AJ+vq8
a3Eh4+jBbQdSP4E2ZO/XTqXCv4d0pRMhlYYXca5N9DDFf5XwWh6le2nSrTAnUAOBK2cU0mDL5XTT
R26+314uwcbrfkxJ7Qhf9uTY0eR5BPqQ71nxszkvkgi8HwUe6Uw6eR0mfrhNvtbSUGCTUJcEB4uV
g9o4SRDAg9WCgMiXyAhzMS429Sv8f1dLqr04jLegL/XM18P0756BTvxFfDkRVH3LM8E0UlW0RP0D
h7rsDHPRhHJFtvY5NlBt26O6XEwlqo6DaAsNeMauabY9idOOPxu2ra1udGlPCta6ZUSK400uRsWa
hXNbMJmKT0CcdH57v31gRP9pc/EemJC8qhhDFvJQR+SgWAmYDDhynM64jbHeod8ZGcpL8/KemJor
ne0nB0063ZXPehix03aSX909Au8ZUSKDeSvTRQvcdq/6ah04eAAgVnLdEnjfJZpsNY0kAda+qQq8
8grxmO4SaFCeHNpE6qFtzfGYJ/g3W54CprEa4LAR421lCKi4N/A+Hmn2mq2onRyTu3DA8938d9Rd
q7yIwDQXqsOonzUiNmcvb8Bg7yuJBuZlP6DDdzhxpYl2U++pPDZWFBMoQytWOc9R4uLwGIzTvLP8
zh3XKvWdwRDld+1F0LnEz5KJIkNPm/NEQ2/FAacEQOsVqumc6X9u1hCxJuHJIgGxIXx3TuWISAuL
RzhYpobdAOWqo8tepb9glSCZEqXCu6FOerd+lWM1VG+q59imZTJaUkQzBIAtjuSfFdq8VmQHT9R7
olrXDDLx96v3yneSiyDtzon0OaKAFyyjQqnkcSBrtPTW3gH5MIqMYuqh4i5jdf2IwlrbJ5o5vjSw
0k53WZ3Jr56G4Irzd4MTcP+7Jf85SU3PbDWnCSMnnXkRXQuKB314hMudSlJYh7kC3oexgSV1IDKl
v/MjXh4xXb3f3Hq6VPtSC5iaRzOIV4+5QZK6U44Rnk7H2gQtIici89iYXf1WDXmvz3TT2wTfJ0uR
647LURYGzMJtNF/PJFa/Dd8p0BOJw9rehBO/MPdz8y6zI+4Om+ZuiRAxT727GsbUmIHO2CHLDq/L
ZHKr2Mw5CZH1RbWdbfgXSWG6WXiN48PK735OdrCKegVQ+HxzwiCrW2oW97Lf/BnPt5ETedFu21LV
7U61tPpdSLr8b7g73WyyXpWRDRTYkstH4g45ZuIIyt2h8K4MuD++POf0hTbqN2yRzqeVXuz6DuHr
2bOPGYRxFBPyjjevE27RSSppxw9VefKj0/48IxUu0VOoLcDeWZs//oH6NLrnPP+a7vkfp/FEu1rM
LLoqE9vRcC5ZZ4wIfSFnsbPKIXKzrn9wOhx828dVHcoAHdPJHwuT/1ZccaPfNgUwKbxF3j2aQm1L
GkXVIMEH0GzW3Yj/xa9c7+SSEjc4dY1yfiDwGYJma93ZIFIa1xJV5Qc7B3o3gOAA1BrGT0VyQfqI
y+aMGI9TWz5syN8stjH3FDucI/SdwJWrc1njEzCIy2O3fJSYOCKwF6n7az2fXDPbU3Ql3bHX+E47
ZFHOw3L4Ollpj8GGsBh8sMGgn/EZ8dxshuTEbQ+zXNenrZZF1wr8NheEJLzIBWyIWFyysy5qBgfy
4AFhYAbZF2DsmN4V+VxaSnQUPC15tgu0GyJr/Y0JKKh0dh7T08JAGqbWGKF4ilGZPKEOzbt7V91K
i/8BL86C3MMOSGKkMtpqBDlRRYFP9wWMeKgpCLgLbW1iUFFBL5vXcvN2Ocz3wVKY8QKuZrLP4Ar3
Tp+jcfu4735LK2AWRAbEv9ro9GkC/3h/Qtk/d9o7Ib/R+pbgXzBi1AgIw7G0xJvdiERUjemr/joW
AYWHDADqapdAIlyvwziDsS/3dxoIrejhD5YL13raFZqwlPkEoNSqL4URcy9I42Ds0QLG0ztm8Y2z
DPIkN75UZdWdBjVks+0TRjCsfkzLKCZgGxjnc7pGuQ5VuqZslVPrvyFI4i08v8sCiFQPNx7kIsoW
+IfEMvglNUQQ4bCm9w65Pxy0HIuavI1zWc9VSzhgMF8LZcYHYANZL9JdJt/pJIODsDHdIJQPXYGd
JXCW0HXHHCS6D8Iwfz0LGOgqMn4LtkOiSeEqsVn534Nq+VXfamq6zgZ5gXrD3nQx8XCsBl9GMErp
VpkWIuvlGqpzmJQokxQqX5l+G9w6bQ7+7yXPt+zfu5o6ZgGLCRDFtkNg8cecGmjIwJzLmDAv5xcK
eOqqMzl/CLFa5nf9Ve2/A1shhzEGiyaT68333JHh7NLUaSrKtOxiP2SzsH+Kh96OXEMtdceGMbTC
6GYfG4bW9vXXO/mI7Js6vD1p+JqCOcZQp0ipvNv1QxpTXWG8lB1P5rs2ujsxdl1qEgUC7UMjkLLE
OxD2yVNIoC3oP2UYcJjnCHytbtIRqAp3TR6/fDnJLsudOTv90ivUurhzuB4yrYaRCDpUovd0YjEc
JgzW4v8xPB9fyD4zXf99mFU1rqBrJAevBsTdLZrOt4Ee4AepF5Z80DmMJYKzP9HGaCg2LjIfbNHr
eZDuJFw1w0W1kU2e+1KB/IlbbacX4iAWpqqq4V4K21KQbOUmjDebrA7qaAD3Ql+EqHk9DkNo9BLd
CfForc3wn9pNjeonc2ZmucamRIbL295xgle59+8TgCKhsMc1taNhBbOlGPGQv4QLPb+Xc27dX3bb
DqSzBsj0jCiGvhdnvv57yc1XFqw2mZoLAidhbH+/V8hZau+3zcu9UjWJiU0pBq/WDG/jFH+3Mx8R
CUIhxsB8PwXaDUYOhYUwMpBIkdsPfAx9XzbiXAAeticC+VFBUqzx1PPz7U+scle/CFG5sz8CsH5i
Kyswp0+t/8LjXQ0rINj1nnsgXqpzn55SzPOC+o8ASPPiZ6U46KatzfMjKI1/IXZkkqGCjLxM6Wg2
sgzlz0UotqGOFk+5kLiM5DtEoTm+bun/GNMSyf3FPgvzw+//ZMz9XYMHsDzXmcg/H8oitQfKO7du
x+L4S7o3TFuM+DRjDFQFymAS+2bXrSYHHPxG77UOvBOxK9JjZJ7opQY8G9pw5RguMQ0Yz7KZLvFB
oyUsJnYQ8+oZ4kg/qesf/7LuyAvT8nQLqYrEQx1M4wmhJvf9DRLrOHn44a4oCbYZILTzhVANxIs6
aJ4SWjJdPR2RZwYcfAgy+pKEihpsQsLTx+tNN9XPXfQ/FCyrAon5m7dqpePzV+wXqE/ykoYjv5Y8
qPTvuX56XgpiFkFSbTUpTrAcfA5NYJOW23NrPNWs1xuR6qHAmdMhOZ/0o9ZExzQMcqX96LLe58dS
uqHAi/dubUmpvY69jvwZIbI8pRRpiUg5DXmf7cPc2f0ezp1W/100qQ4Arnanju/j89EYcefle1TI
fnMmyhvH79WqoPpaN0+v3lQ430XkBlHW1OkTs9/WxzGSPjKtEm8CEXtJxmP8iAcUVUPzAYTcdFw9
U2PsW3zHOeNIXsP9rsY8kEjtEGGGZzshR2jUSM09D30daymmumFD6fF1K6jHPLISaTEKiOhzvVcI
hO0fDxJ2v9M50n+6A/O1ZM0WvdnV/fv1FZ6XQJ2eFa1vca3O3ELhL8U7R+RTUMp68OrtyudBcyKE
8R534GBCfk/7N2nUeeHoLvqqtkCthyXp0Rp6/MkcVr7dsWS6l8Yk7HJE0oCC0jKjkad6xL0QUHK9
6dx3LJIX0SPYVxxw0/Nw0sZGbYngung3I34y/zDjdUPPYEuuN25s/Lrpmgvov/MfBRLyZAXGrumi
Ti+lWIm3olzqbVl+MAhntW8bwcczZ34YbfFityNgOpNpwif9G1q0LfzyaUFsiQfBojg8VegKx/y/
4DzXcaEQG2/accUvpOukj6bCI4C7WDa7miDOBRoswi3Hm4Vvm24IgC/1D0Gl1OB5KVOFVrAwOE0I
m8Kx4vt9gjqQ3S2jhEth1yMwDvQfMmZTIg6ATjJX/8yM/4bOyqtu8Orb50rfQcyypArjSDuFNgHy
dQDLE8WWU2JY7VsriM1ADyNsf1taYyugeB7MS3V4KBeb3bMLH1jCkrA2qRE3nyVSBO9n1Yao68v3
cQ2i/ErFfdOK5MRbqNySyi1qClqOwHj1SN/YQS64q8PY49BeHeiui9Q84y/ytwGbtIC1XtSMnscR
5SZqMC3fbMxsQf2oy7s7WoH4iGEPNPMFocXLyYuUC74rqmrnIXfXQWetG1SSfvVxnnUoypnF26RJ
Zdi5DxHqF84VrhzvbzdF69kb8OyXDOfr+NWk8GviRQCR6VN2Z9pJ45PZ91pZaMWMEGVXb+g6cvAx
fvAZiQI9wjjk1JTxBclFeqJswEh1hgNuf93cANZ0rUJl0dMC/SVP6VIuuvQuUjGTfU4VH5dGWl3K
VBoMKh2C3D8H5FjCHi41/fK3k3pGzjHfr+yl1YcCffAshTel0qVr+9OgegNVmrPhkd+ssZrWL4Yf
VZcUbKgVpITW84E657kTFJo8FRvPfCx5iTvyXVo4cO/uYENov9rHCxDZBaidjvt5NAA1rzUVWmmK
mW4qjRSiQ7SlFwXK/lYPQM2XXcA4uyZet50ZSb9GAJFswcAY1lv2PtfY+e3j2xQ6fk48dOFoz+x3
W6ymdJLbxp3F93qvWuB2dPwbd+MFuJUeii/jEvgo9SIVWqtXQIBLzFyU8uQkK7AI/rpYTWqEljdY
0ZddaZsuf+zNytS0ktXOeUmOVAUqrUPgIJ/AVIdK9s4raHj+EcWEHk/PC3uDt1XnL9nHF+1Yb3wH
boN24tun0uoMgeJIO4J+8jUFJ9uOKUQScq8F5YK9pAGefstLomsE0bP8EIqACKxzaAuHBYgBqOWB
qCBApxt7FAebyNdk7cL2rZf3CtBsQXw3qCWaWXgjItqBPy5LjdOh7N+nmopRiXZgY8yUBe6aWM+M
HJ1/+cDGti2fo0PMoeBXGD09eIAj8QhcR94yK6tzhE3wObelWn7FSXV4MJawJuPiO5jz9C3THSaK
xbFtKt8HvBuRWPoZWRk5VmgATNtEKQe+5effLa/BwDosN++4HNjb4ow/y8AtiFYgx3m9OB/gu/Vl
Po4KG2RkXGIFgtaXU62ZQ88ArnhUNIElTVK3NFxqkJIUocNFRqUu6IC0ertfRvjQkO6pHhjV7w7I
NMTZnbYAPRE8aX4veKHvzPOcB1UWM8UR37N5QgxCqD79kMrVvo78mIpwseIpm9xQokKiUIbC2UqD
SoR/XcUKBy/GBz67uNKNB3wiM/cxVSheMxBDSLUsU6IIssgyQx5Cc0H0/LBaBc1u3b1/2zKs4hgR
iMGRH9aqPvJbz376S7GJaM0Ae3oX35V4Ck2WrR66QV3ExJhCCL/9n6R7DM7U4kRD5UOQMnv7rUmt
FiEcdnRvpXIP/a4xfiwhTsAW7NoZghkt1+q6w7zEnpQtuzWA9FKSP4xFi7LLbHSpZndiwq3/corE
nfHPwa3C2VLwYPdjBtfNjWCJvjccHSGPH7CEKcOWzKaTRCX0uUVjBrE2XFcCfRkXfl+xv5eS4cho
lsNCcXAGCVJjh5MB6bvd7pOHu+fuiDmXqjngM5RqPOo/sT3NKo2zS8K52z3I3HlM3wsO17VRPgJp
xEiRFHhhQaEb8RAjWI+cGWoawfKxGtAum1WPNNjx89ClYevJav4JPm/+LDhu1K4i6u+7KJGT/9Jz
ZgNy8MKLENpfGeK/OIYD0d8c7a6gvwKHe7rlOrOA73GG1FrkYeSNLK9NqQQD+Z8wX0/vn8fUeo/d
bzxLXW6SrPBfD1JZS7GTX3EbFTOJmusR3QnPs99+eLsD5jFVyr0SJWq3X802MYmnp4TZcNh5Bewi
drbyzOS9tt1MNVb7sZOq5UrItGBV5Q/7iaERdro5sw2hm3u8eRkcMJUyDgAAxhgjl/VZXQXIqBnz
Hp8MgzbyHfyvIP9LeyEkJWAWcm0L+NE8SA8zsZuTxoUpy3w1eqz3yjQKhMkB7iwG58JYXy4DqmQR
s3vUSK1pjyScf+y53lWYlhPd6Jk6ABmKVmfW9QbWRH/rwreMYns4nZBD7U/XnG8h6wXqGznbL6PE
SQXaVFXfyawxvqSrgbogY5tnM200hDn13wYB3qw4b0udFsB/JDBxgnx5gUIdNG04+uicRgPNQPY6
0tQlq3UJqDm+/EtCfpzHN4ksZFjCOS0XYPdUj6L/O/cCMAdQWsbT0+DnjI9wT8Y1pokibzktDRBH
Ihczqhyv7RG5ffwpvjVynykQrq21OA+hmlH4wPIrW1hc71uhkV/tEg5L+8KDmJ+cpl01K7oZzHXQ
GsjjMjZDCqC/JpP7c7kYgcBpagOO1QJsKkPUY3E9p+rNGc/ZKOK7ngLw91pPIFZcsYJlXeIr/Xli
YrO10Vv4Z1GpfuPE9a6TQLyjQeQ+bHwQB+TwV4PW8S07Y/AH743gb0ln85ziAGwBE6Z3oHLZmcGr
BVD0auhO0CSl7MZvxKC14ltX1fXTKEkpXs5hEIpGXrLO9qNWGmo0+CjXzfhc+sbaTcDF9C5dOuIx
+2eYmpf2YDGbi/Ws/dpmxIHs8odgLS6CtGwXA3RSxB0HujcdVNh9YQ99N6hXEA4EwXSNq83Mmim0
4pC5WGVVMfr4UdhaSkkH88IvBcEIwG8PdDymsmk9tafsd1hiDIRh7SVsQsOp1auy48dGKixBNjas
sF5el3lylywZcqtq77JdKop77lI1cpH8MFyjuNuiKxMvnRRIwDQ1ImtmBxj6C1UlPiw7pdRfRVu3
WaVE+UcGOjxVmooKR6ATX/younGIVOOKhxcwpQDPNpLh81np8H60QEOZvZwSjwhnoKUUf6Ih38Cq
qFhGJGve8afZd18UpJBJUt2N9A5kgOKTZULlU3chZMUB3nxm24W+TeWkuECz2Sk3TWed4jWAGtJp
N8v6SCM73bSdOZ8qklkD7EkaAFzzan3hU7QzdXfffdB5u5NiQXQCPVwA5YAwK/pKJ6THwfpUIVr8
qFdlSxMfVN86T4CnLk4JZJGMTlTHuvUYgD9kK6e7XqutS/xXUW96OBK0nnPhIXdvFm04cgydThxB
F/KbK5exhOKwFZZcXWgQW8GKgjRUgFwpIvbJ6q1YUbRIEnD/erNC2aaH4KmnNoHvEWGj5fRyEpuw
DWByBJxl818fSWy1vibowIIbcJbZKr/QIP47G0qblNQlUbBYbV4AigQwzGJtCjUWjRG+nDH2fecs
xLhgCmFHaSkOGIEdo5vcUxbDZAHb+pttFdwUrvUiuaymkSPfzeM0xgeUGHzoPXtXIR2EeuUwwAlT
7f3jvFSS80SMAibyNxOfKR27U0kx1WrJ/dJkpwSt7hBV6eq79SrT/AmSBIYD6blYCXfAXmMvUCsl
7mGITpZJRGmZaiVDw8rBFIb5ke4qQxjw08YKEAxaHo9kfxPyGjJNlSCLnvChaPbx357fUAaDzgiu
zX8n8EoT1aMl9X0MoZAl5TTBTcvqNiMgfjY3Y9FddhI/fsKLEDZrUrWl8XyTbjGEcpnJyG4ouZ5P
1TQYaBTh08a0UrWuijr4ZrHOcUIb4v+I7F2BLvQXzJDFJOK0oBwBtbHZ7ynkw/c/4/E1ShNjDllz
RPOdOsKotPFwv6/2YlO8k9mYHUNitEE9+xE9hmF6lxkafKDZU2uoQ663bQLnIQpIwxHicZInhz5p
ObiXVSMK2rznvqWMWIOSac8G3xHpEqmVZiiosfqyD8JSdSUUKHsoqrJhYx7C8gc9sixBFdCdultL
CKsVzCoDEjsNTxUquQxJZZ5QgXr3Bv3Sm8Z9yKfiIu5MwizCTXE3pdF6x+XU6WRPwxTe7y+MSod+
IJlA2qyFo3bDAW3tsiTy8MyrC7RjorzhCmpC1IR/bBo+I0HtVnre2xjKvku5iXYG9dJ2difYTG24
uNLeI/cS9Jert78cGGwYu4kVMaxQr8C/LPDkLJJGaYpsYAeoasFZspqARATh7N8RjLpH7vLFMWx9
YWgWG3NZf7nJznRvcBO9QElEDVDYdrnyPGXErYeLMp3eTI5u7d79bNzFQYzmlJbpvIaw1Nhaqw2O
eNZHRFBXHb/tTo9ognsgwXj7rNC42ihdPe6Gwjn7J4zY46p3DyKtfHjw0FHPjEf0uqTCpFeWOZ0d
/qkOnsyAXdNcc2LScE4raFj+3jmZgeUQ9x1yVU5BDzbOloh7YHxuv+JS+AiYO5XlB5yXK0CMKq6L
4FKA4gF1qpbr42ewWpWVRxzr0LzYWklkW302BLyS2kQ5C5UGdN6snnS+d2+K5MLboiVMIjpGH4/2
Eo3IVPz1ZhiWXaN9Wnx+yB/0ZHmvTZwIUKLPC/FeADvUOw7Nz0cHGbSqMzHMZdgtaIOzrayIAicC
pFHJSiEHYkcSIpcMHFdfQk8PE8ydpiAZH9ifXwQ3O3GS72Sbcp4Z5AJvFlygU/9APdHT32UAAIK+
BfbnNl4c8XvmTTmKe36jP8Ya99KEjuIZyRLZ0EYeIXRsqMOtxh4NRlOHORD3cQP/fdmD46J6qlq3
/hIzUtkrKvT/1F0EPU6rjLEs1sEfvz3Rq7BZKy1bb+eWS1X/pTVZCzoFcI6dnhNip1LjXAkmSFf7
ezPWWZ2Pr9ZovaVe2qKNkumLqn+AmcMLY3oyPcOEU/JkwOhEuLPq4TJF/adY2i3fiv97xwjmjIDf
M8Nc0Ueplzc1w6ZZtAbb3ASjBurla720GYS3ODnKNyf4vB8WTWUDWSl6HhGb49rkyO6SXAcezuY3
Xyar5lYbks33+FJWmkr48hnjK+03uqMQ8SihdAcBhyS1bBqSOL7/B/FZTCzuRqWTa6jMEo7dOIeb
XAVhWLAjD7FIPsBFOtoLtPWAaJdvwgV15c0QzOQ7sKU5+gHdChFt/3AXmMnfneaTBZP2sMHSwD3Y
6K9kgxuSgxZsL912RRS+SbvrMaRpyiZdbDFBbRUBOcUCTmS5Rac6DReks2gxWABdz1KDAouEC9op
22DFmj0MtWprihlaSJhyoIrdAEsKUB6EXm3P60/6yKc5ZO+x/w2r4eeE1hjF56qFtM5hV/Zmczx0
6FEvAkgTsRLLMQKniu3Ptj1ppePtvozvkpPF5Zbuv/cQq8EBzkyhHr4xOWROdcs9xotgZQAtKy48
7n9a6V03mYqq5lXFvDEktKu9iL7l5Aj6+VfqkLBNuLApiLD79eN1kK4wLDFORpHmHFmRpZMnChgy
lINzBcQnguq0yCshIhkUPqyTUVwXjNF5XINQO0Meyc2V3yF+5gKDMxAzdFieOpXTnJmwQWj36xCI
b9yC2AdiFf73i2eQOXQFi6gPPxC2lTn7JoUSBOc3gtZotXArIYgr8Vmg5syTKvDP/FpB9hBxmMNZ
HMjBfAqVddoMP5TC548ExQmP/vpA8AbVmMDpp+zLlfpQfzz8ctLb7u0zZAKCngAmyqaGi8CP6UX3
6ld08sa+dq4YHQhB6omdNzbcjwGdEEAYXtwxUZdWORFbI1/JTQ0QZvx+2hkuLgX2DMNCAPoJxhGu
AXXDIwPOxsOIO+nPfrAkBj9bcNXLkNVYZ3tDvXIFKhipB+zRygQkYWKdcF2OEFe2/hIQ0A4SN011
GgCwSzjpnLmPGaAAsJ/KVJrPbzlkvOAMAuG7MGBfb3VBCnXSQuPlFroaQWERG3z/V9UPZbOgon7A
fau9P8nK/G+Mmqix8YP1L0aagK9Hu570Ncweesyrd/Fm8kNnTltjc2U/AtnyeTYww8ozxlijgWdy
4TxBHXrzo9VEbeZCjzTr0Q0ZadjvbN3ttqrJXswmToX2ABFxubujT/QIQcMgiRT9ghsiv1ksxyYb
K8Jxs9+1ZFk5kTw9S1xCQYdmAZCXaojqQaKlc1JF+itMaHJkfg3ev1aRuENXXPwVkn2xG/c6W3ks
s0v7xw6J0QbM7/snnCESyaaaD9o9BoqC+wNfYEK9RS6bcqSTd8+NSEfP3GZE3+0aQUPrSgcSugD0
jOSJZ8xNqqOmCrKyF7HqdZ4oRkQTZzA1jzRj+e8rE4FlgXJG1rV4zuIdYzNWVnNi/bHkyzhU8bGs
GCB/B6FnQt8Mr8vIKmdgX7heimV+EuuW5VVf43cC79CQbWHWHFG5PlfnWcWQg+go0jjtfMCTeY5T
G8f2771ySSl9MeWbJa+Y50tV2drPWUQwBnr9emj2lGWBWMZcjxsn4RPpHNyuvaqkd1kVb1Vlf2N2
fXrC4/LfW7N6+u+H8Bj8wpj+nFPN8AB99DvWq6qWh2DrBxWvZALWtrlIGEGeGg7RpCfqWfHRy5ji
2vU1puhfEqsqk6f3D+HRmEzWQ5UtDouZT5awapc38ce7JVTDDJ8H4iuVIkOMBTp1ZrufBio4uOgc
/EqK1Dukyh73q0SyS7yyyxagqsJt2Awk9J2Ujzd6ZZQ853ftLa/9g9u6zXE7higwE+rmVrI2LEkR
gAHL1bQJM7vIIMoVXD0CrKp4JqzwTfpYuRtq22epz9rjZRMPkf0K4FDmA9TZwcQDwEuvGdTNQIJW
TMqRmRZvuKRWVaJa4M3h01yhhv8EivUS7w994dhAxJuZCd7FLmCptR5oSM6yy31fhOTikIHibZWd
S39LzBN6Z8gUPLSVlL24NXM7I4LvP2ZorzqhNatDh4fowHIf35fGp5qbO2Ym6y22+L5ap2dWQrK/
5I+pS3x7426kUcuJxAqt5li4psSU4mr1zsUethlRq3UTZLyGu0unF7aU5kYZqogWB+I22+V0bZxg
yqXsGt2s51178lXd0i6o9xDkrbWOrdJ3KffenOMEJFXWJzKXJ/ik4IC345Y3YbO6uO8/MiV3YTLy
pqFq8YLArg5GP0LNAuQ3N29zb4UtW58AjS9VjTha2D/zf/mIWiW3zHUKDU9vVK3yBGeN36cHO14k
rgSrzIPFZpwzlQOpgEtAh3J3tPbQijcJ0L5MNwq0q7rRaqbWgqyUTSCR2iBwuYKOwdU+aXHcT+ED
yhfQgj+TzWo7JyLC6L7NzFER6xLquLrPrhGJOQyvyDTfFdxZXvSMOGyMEWZs9TXPlX3RtJg1VkSl
oMtuv9Y4uNBLIMYZOErg0JrccTAvKcQZesby4uNJEj2aTLf1ZV2661SxRbE2ueg01vaSrSoxare7
9pASDSiwlWkVU5P0v+BzE5U0iIJ45ua1hz3GcJJTfBn+2Yi06GEG+tH3ng5FnsbPpjc968eMi3kI
xvrW2mo9DTZJ2RiS9kUDbamgxwj39zDy3F8vj9zhgelrOtqSsSS+eDgBJlev8L6SGM2TkS9eizFx
GYI0/sWM9Hm6W+RtxAjJUGr1w+aDQv/RZ9CsG1I4WJrZhq3TgzFBzZit9L7aM4Bx6Ym3eekVWZ8z
WaZc4/U8fPx0NouIwbw6VtIOuownCsQEDewlIFpPfcBUiIdzf/uSDCroKAjHDICWYwRb7XZv09lh
ttypPMHIR8Gt2jo3q2Dixpd3HmQm48FewjTfEmQOKTy5NqBtXt9Ea8sDy5tZKobgea3du02VMumx
23OTtrLpiI71bMR3aVWDLhafkXxzuNmrFmiSsNE4cwSkaF1ZwmHORPk/Yk1gP149MTnPDPMML+uf
R7LTp8ZpBKo8moZDv9lliymTC0wRSpHnQ78vysuI3YZPssuaWI/phnANaclOi9VRYS+HVAzyS2Y5
aiep/UfWr/kAICYWAvS+lXrANb++r9nVEVQb7sbVLjUCeqALrl1smxEu6R/7BUewjCfdCUvlsTqN
VzqhJTo3AvN5X/UyKiUqlamCNZV99sL99vfNYu7CaGTrzHdyYsL0UHuI6BCORrsFN40cb04R3d5K
vAFKicLfw53zuY1HvlZyQaEp6Xomij/JQD+1jwXb0OgxQuGReaaN8Agol2fG1ZgljstyK+neUUrY
SBYwnErS/SWI+Y0GVpLDvgIVh8rwtt98NVtP38lrb+NvSSAGsU0pli75eN9QCFqYb2A8GKz0IcAd
U7kIWBuMA8ZfZ86hwS2UwwRFRVEgE40uLwcH6Glz1iqJXB2oalteMMDPtui8ZHP48WH4xocwOnGQ
DaAd4UJqAMygueEwDmXIgE6JH1jwQQUd+1yebYpADsD0iKM4tGrAywR+CNxKcqnoN5+Ef95QQLUZ
YtouLh80YapnZawWz54ubHFgKSbhezNTtiSdBE8U3ciourS2aRaRvzm4HOl76fQCaaQZXpOXuGH8
5zlP+8kbw8hG5VPHlpKM2YmcigRHic8LwMFsgtRJ4Sf941jcBbkyP8rrtIiUHgwkH56auvrwlLey
evGLsAk2TNbRTu/3wZg3h0lr5DvCsaC77hfVoZw3mIzZ05+40Hz/cLTvb0u3LEA68+iht6k4DwEB
CHfqMA2c6f6RfQBqLxmczdIhd0XVFwb4LiY/yW+iXAW7kBZit2Mxe+IAOdqU26cKsxpIGzLTemTN
70S3QxsIyQgX0DXPKqTrFmoSTozRGHZd3m1SEd8dY4plBzxZXiAgqNB6Gav0UYL0e1ZsvTJfSV8A
rtQpCgNrwhca0+/JogG1uffXSfnhEC8eGM5fSAjqABpHZlxDYB4NzFtHkTbc5SftqtpfFZi78orV
J6drFzke1IBZD8DUh9Bf1WR5pG60b/8fik0gIJCg4/o8FpDq6HM9mez59bn2NekGi7XuvRof4rfC
KxZwh3BpW7dDPjv5VHT7GCjWjTJ/8sNOFYG2LS0m4/61XQJVMCh2WMP6yKEq1IXWlNUyqJb+ttic
FMdXSOdrG+nxhp2N3EcF3P4jdeTWg8M7rbWKhpZ48XjdRHv9JOVR9JanOp++oC2o78sG9eog0fMr
HrFG/U11NTdrtN6xaYWGik3B8ZMiyhXED4Dj7nYBLQcAWv/3HwehtI9As21Ux/yGpLJkciwmfazn
9oK9bbGK+t7q66D0u0u3veVoGdFLM54U1YcascYCYmA+6g9/hUj1t1ei9oxdnBsftTdreZ0837LU
EAsW6h5MFw5rjat8Nr11lKyQ6ak3AMb9xhRaSI3LuLOavYv09F1ie0czJ2ie6xTa+k2waCpnNbWx
dC282A2L3KYJrN8DIVysCj+/zQA5Nes2D2RBAlm1oxw72jK+V869wM1kh0FKe4yRysDfEc99HYn2
sP0ur5aOV2paXVzfhuE9fhJx2KpSZ+k2d4HZPJxFbibaM1rz29xyJWS5++ZhBPObuHVM8b240ssB
TNkDxV7HuYiXsyRP4HHIvwKeKJLSDIQi+b705tmDhk3rmmJShaj6OriJLbcqEkB44VPl1wmpBUTl
ZUBjhlXTTGeC+wzFJD7pgs/0AutY7FiFLKr2+nimgcotL1UNjTJCWzGbHuqC4UmYZCzMzCehH26E
lf0UnEJb6Uz6fToCMh+iyQIAaMjkpSA5sYnF1bEDq2pq1jYaFhAjRCTtSrW4kHonqfVWOv6Q6Xn0
FVhxNirboj4FsmU2L3Tkn6Hd1G6/qSCCvEEIMNbigAsQgGcLGH0Oqmrp8OpqE4LPC9VA/FrXf877
xcNAGBNzHo1u5v6qm7Cvu/FWYfKxEGdqVJhaZDuQ2jMvSDsRAdZhk1rJmbVEGtlxUXRIh+OzBaaj
CSHhil3mHyy8ttlPm1WgnhsOGR9c2kjFgWvooKvJyGvQVkx1KMMPAslIkYmX3nhpiMJvJDNY82C4
nZJS12M/qvvW1Z3MKhO/wHhHxGiPH2t78zO9q0bTVQQMgTvl8kl2dpByRxmRx/ruB+E/amYKkE4h
pydlzG2CZjVdmJhyzcXyymZvo/wLgWrjo7Hco5CeYfd1oR+zZvjHuJ8q3CespE08AMg+CpS27U3S
Sj/sT7lIntd0jsCRFXq93FIxfQlqOnzucYZpR6fWQ8iAXaUZFjymLDes6tZzeYQw6ukLaMRqlWiu
5H/MIWFDgElGBNC0LENOV0LLWObOs7dKZgz0l/3YSAtuTkdooo+i53+y2AyjAsSNOlAr3MRwmuGu
zC7Q8XL/zS+o1fWa7Dxk9WlPNKD1VZT6/X6u2s9zJWJ9xKqCPO3Iji0Htci46KVdTSqgNrKinVlp
vnoCUrmM8k3fms5DoXrvg/6ElPifhfkJFBp0t9D22OxY7bLXdDyFCDvDOBo0AQQEzEqwxXNAI4Vo
F3Pr79iEqzxXNKWpCPkvGIIUl89O9FqjzU7OMeKvC6iD8sh12DfzGruexZwyOVEwSIC/z70Y76AT
Bb73FOirKRTQpg/LTDRgY3CjTKAuiTuvsQErSNfHt05tsLg/1Mkx16w6ssVbizR68sc8eyMsn3nS
/Hs7ilY5WG/MI5AONZ532wfXGgCoWrXgiL7Vh8qnkkjqZzwgK8t2JosRBly9R+ZYmuajavazbhj6
3qLG4S3tFa9ZoEGL23JMN01/KEbsPLcax5zr2qM6C/OAXKtjcMimwC6BKUnup+vDz+6HXDnsQ+Jw
HDKaZ8cdcUChtpzAJylGQDSsitVbjuSERkDHZNbsf605LWE475iZl7XtT/18SDXadOnKlSIiTeuC
um+6TbrOPUTtdqyz0aPcFxxiPjnf5ZLzqmFNo5dNm6GazPvvClPbiN7vmHfw5nxiq7t1fGY3/4pX
AN57L54elNkCCRrEHMPpPqtG8QtA/GJ4rsmYsToGJ/kr9kdEmPB2m9sAxXmYrLMnJeqrh1+s/N4n
rF8SZKhgt7I8NC0LhnUukMzkZa+FAUgXROkFpDHmXNnTmX08TUDNp5HjxreLlxuq3GBCuaRH8qC9
TOSU99GoYyT9xHBhV0pO3qu6RFTZtXsmsuVuh/xNGDL71ffpSv7+Ot95UU58yhdSEC5AyXXlY9AR
zvfN8wJ/bwxISVzsu5O3okGVQtRAUxw6KiRkH5Mj75huCHzdXIyA8kBgHrMD7BoNgx2tvHhnb3uW
n2xNIaVfqy4HbOZbqaF6SogfxuHtesh8W8Dr+cxhpp7RUy8DUwKQNVryFfMlON+cW0hiRAJ8QCgx
hfq0iRsPYaW922u2iJ44OfIOBC7Ag5OWmrbP01W8zbvWv5SyRRsK3o8NZD9d9rN1hoOja4pW5FCB
bPOVozUdBfeiEs8ATo3t3pP41xvBkU3KC7hRYyVRebNjqgIar01f2bhWcfEAK/XSgLuS7H/YuKbW
dD0LTfNSeg+r31t0nlOzWBSkQeAWUg7gE6zMjX/VNOCy+t3RdH7GSI1GMv7Cm2gfOHdI3igwCQqw
gdz8SP4y56oXGPinmlcMeu7AaezJgdkP2v8idPV+7dlhstGdQH+sQlF7hFDdoWQNyr46qdsJAp47
h5YfQbSbKdVzxOxyqag4y57UKB+dUXxPW3XVFOm3E3Xu8MjyHwjo76R6Zka4IUaV/VVb3a7T+7Bb
6NPWsGZ/9aTkA9Z3N9rRzYRXLeJdyelf+3s3QvTI8RNHfDToZOswWvdpDH3WPzUXUYkNNfxJjn57
bi8O7xvs3VxuN4E9S/3NktkNKCBRBvhO/twmmgq48egyoXL8VFygD38j5vLEJ//IdEErIbeKMG67
pzDRYygqwUx6gE9oEjl7PAddMNy+enGM7yHKeF8/TCHr3Kj/DzXFILmC7rhj4fg7wKohNpl/vmBe
cesBCDlAlFZVErfB+0TAsKLwTCxhup+/S7c2mbBdxWty3hO/0BvfWOiHAZoeELeNmIdYMT9FPXlE
EaZXEBJJmOsTFNuACXT5drIHYYmBcl74eqgROF+lJOs7Yi/FyOCALUMi9cQZem+TG/GlMnJwflpM
4ga80jySAbc587O3hNWc5DpIunKrn2W38iT6CrCLpgdbeMtWUq1VUNzGaJGUscGj0a5qF7hIGgn/
BMDEJj0aEUjs9bgrH9tmNzytoZVXgrn1w328FDmomZIQbMdb0Xopg/ISosiYYh+g/bCkayKW34cU
38zrR9MmqvoI9IZ227zvGwjOVVv0pNrXFCXm6xunmHDeD1+0z0HKBcTwQGd/Qre7cwggCrJwGI7a
JST2LDXOYrw38yk/K/aeD7tlkmupGqikXe6WW5yGmOjDn3QNaU32DTjFTQBIzS2BA4xk7KP37Whp
MkjYQAFrKRGaeE0cT/EQQnE3UzOOn8GC+3T41tcTvh2gJ0MCFdgcIoHfOlzNktkkppYREcDVwXR9
8rU5HVeLl94tL049064Pu1vXwTspSFcxpUHeJW4HhqeC3Xm33nCpOR09juzXPd+MQxVtaCm0cw+9
7MvIHrUCaPMVvnO8Fke/r5hdKJxN/R8ed4zxsTJKkZ1l560HQIQI9zuA/ZgJHuoz1NWzk8imXUoD
o1NipD/iMsL7DjTK2BWwXbzr+n2ssXLwma889IHFHGQE+b9emAMSxlWwPJO/7n3z8YQbEosfqJSQ
shyqHsLacPecMglit2WC60fnMf0DEEcRlWfblZs2IlSOBM+U6zgHLixIKP+wBMqUgFhZdV4wFrrY
5tEZfcPzqkz4qkD3pMTWJOcLT5aPPfi2ofc7q94rDDIukpyFBsOyj5GsIvgsI98p/0VK1sp0tAh6
9+pc0QMcY8cMkSzY7+MTSlFwUwgmUM5q5ZZuife45BdJ7F0fExi5kFDii1kNtiwQbNXsJOZaZbEi
Ih/Th02n23y/MyFiMAOI6Xz6k1mx2gGDZDxt8TUS3HH7MEw+DZw2rEBqb4gHMgM+IdcgXKhhIwm9
SuZqV3lAz462D4tR9v5uX1/5uCS5WGC0bGZqhD/eABMgXhFqLj7/nDGgkV8YNXWXN2sauZRip2zE
RGkx5Nb2eXk8WSu7RjpzTCCb312r+kRGvWMnKvj2fz6WZuthkBpNHnntLh6llOzyMNzT9gDjkJDt
esH3HPIyrxYvOg4wTA2ySk+UaDXnAlfWbdC5i4wygpHxaOK4kWWIPmgMXTctNaUXoIiGdtKQBBgY
+fRxSYHO+iE6gVuMovjOiB/D3QBWNZ7Fp8nB4xKwOKUgfAqKnJX3sIWt5mBcBvhS15tFIzP3xdH4
rbzPGi4bCLGwQQkAO0vmjnlu0uG/7fAnzwlUGqLQVQZzXxlbfY81eOKLU2P4Rjhgdsi6uQAZDIld
6hx4pWhQkG6HS5MZCsHkZZiD5zezmWO0qEN6s/CTe6NZJs42Qx6ICz2L7hwO1c94sGd3HHl6pGdw
uAqeGdhStFJSoKwAf24jNE5My2h99ekmG396vPAxQVmA7qs7tQknZ/CQbRAzFCZTUKzRTxDg4i4U
iZsAoTXxPSNFmINqR6xznzzEoAWRPHelGuJ5g/6FrN7XRAvDc/pGQHvrjrQ2kBHwqFsMXf9Kce81
wx6Emlc0o9xbzHZBhVV86ki6suDqkoxUQNhPC5rqCt6Cuj/fdwdAEVNPGAY7aU108N7RSrw453Fa
Thqf2mp5XDR77ppjgRZbnUUGnE0Wu8fiuEYwlkTPggPXFWtRjTFOKfiz2SNAVO5WufeN5vUJv1MZ
2Pkme17d3nwECRvLoXkpIZNhW78ts0BGGtfMyDkcoHC4Fsyn2r9sCW9bt9UiiIgkEpllspvM9+Ja
OzRQdKSI4gRcrFKps5uuFudGBw4/VKnf0mlCxn+LnWNaTJrTqlaH2RbepZS8VccAFGD9CEsjQR+3
w6lLDr7QtDhv7AjfmFvpxR1/2jSuO1S58jT2qRIXA9TURGDXCUEzU3yiwbfeMzMJjMqXx1FdDI10
wgTtkx9xyDCi8x5tCIs08epd+IGMkGz5MwpDmWlzprgNua8ROn7xA2+tjTNLEjxUMRcR541JnHtA
dnD2dR4gt5fHJ1x9rdRgrkggBCFt7Redh6AOqp8hpxvm90HLbyoe1Xnd/VmTYVoMUQ/jVWJOOIs6
1hpDjVUqKrGU1iBnV0g6ABQRONATZwgJnTEzM2iTyfe4l2mCQn5q0bvpAnnnrchha7L09N+is+O5
qwebOxfEW2MOPSPFxQsEWW2QhKmf6Of77yq4AucANlyBJwyMS5Asd1KCyMwnHZ10Vl/xS1srOiPh
YoBPZNloEjRNqXkdk+IXRqMOfefae994Xmr24nHWxVGdJf0s7FxZEuJ1tHlAVnNmjZjN/t6BWzpy
NjSzDh5NXgTKco0i3netj7Peds20Ld0cTPH6yCUiTFPMgZaFtTqtQldfnMdKRfFKaw7mqYS8hZuW
xVqIDHRPpzCN8jd21q2cw0gD7o7DRvlqDixRtRUGOfb6Ng/dfpwC9x8H8oJX0LHYH/uDWqqeqLiH
VUcP9uZatQbIJenhGjNbVgeSV5dH7b8hpNoyJ2wWzSEhHNn8MHRYI/joTACtVOtTuy4EyiTMjYcM
EFijj6wqDpEqONFGbW9vU+Dyzd/VkkMlo3guKH5ZbQWN6YbysHepPE3BaioWBUCI9p7UpUOhvpbM
bqcjT+nXRCgjyYhpkQZyMIQ53omSma7QYGcs0uU8Yms32o45W8uL9JyvQzhTQzpO9avzc4bl9GSM
6srC6UlbRFPf5R0ejb6y3CiwjUdOQkGpwQwVbcMVT53C7aR+UnHk6Su/rkQN8kAhoivRMTxkgxMa
XtTiQHK/g2g7xxO/LEx+xzlRGkrSD8wwLiABzKr0VqlrJ+rojfQoSsgStMmKLTyLDiQGjPvPRU0K
lDMaRGMf92pLExT2wQxzTFwOhrsp3h3anONT3oMdo0opc3AwC30DbrjJ4QgYQFqa+VFtjnZzay+1
5NKDLlxA3ZSJz6zUKgsfThi2MNU4/OMvJjCw1hZrb1Yp1pq83DmXUWMc3ZxwJunNhb9Pv6LChznV
Rlh8yrbLuirNG5YIHfRiGBXDpPUg0H4gIPOhqhFiWtaBtAqQvGOC0bqyJr++/iUxNuSB1c13lq9v
tdlr984mzl+nHFyoAxGLwW0tZQq9R1Xdbg+qtZ2qQ9/Z06cqDOAR3Saz3Kt1F4nKLbB0gxmHgkLL
/XwkYAfo6ZDa7u5NSEIvlg3OQXzTSVZ96XX44Feu8iWKcY/lf7PL6/4BSsuuw0swS83OfY/vzagT
X4VcioxEYt0IaKUadzULzlZW6o0dTXPTwcYVRMKECL+8GTtcCzdA/fpGnlpxV/I37PzlhOM59zOu
6zhOpOKdQCVm9+/T+2544x//SrhC8CNS5CXJwhPtViu2+wh5sEBFqKiUmurgkSUG20abl77t2kKo
1P5oMdIc8uYZ5aYgRZqaKdLC2FnCnA7FP4oHj+npkAQ5xDKLrUT9w7brK5HUc7AQPRXnpzGgNKh4
ZO2vRKQJuWFHujLJ/XfLQe21kmbXm7nerD2ulPE1yfw9MDL4tQLUHszc3AZgXiwPwaazIvPU8Jua
ekBIX2Z/mw+wjEbQwrIWc9Wij/8W5DZwIyc4+kwtmlTaZbwYXQqjsTLWsrFaxptEJ1ZZso5IfTpu
TEmqmY9Rdj1hXg4TT2sdPL2wj6NGA2YCLKXmkzBzXOjfeLaEk6ScXLVzN1/hEaNhFxX8SMTt81eO
pjA+zBZTWv6sESwHrT2yseV2ZsjJ1U2aTUnIZyRJrtxM7pYUHR9g1+4QsFSXiMQvonGWAzdhlhnn
Q3Bc3sGq3L90a6qHyZ/o99OwOetEzEib6wr1LYGH/JKszjG22PmuL6kAjdwq1jt9ZHuc7xuYuEpZ
9iqIsIr5V6MSDtuwgI1zCPYemHnGGurvktcUZaKO1BV4twcD/y8suJGaLSzh76hcon9id/oZXwZl
41+iX9In7vCuq+Gys6lU+G25ABg4OqGHcUeoKTTH+JMHD6CSPJd7gQ578mNAK3dkpmaT4CYCR97r
HIHclzjg9oXOlQJSDHNSsR/0ljtqKRQ5/KuBwOng79m09RVS0GW8ltLXVmfC3Xwf3KYCdtnPD21e
QdLnCXUalnbBdl/ooRgoDB3M1DXbPTcn1rVB3pcORzpQtzaxv4WGgNutpMVodRPvfG+B17gOTu9g
xFvWS8AQybhOVaXlFg+e8B4GLEQtjj9ceqYMNPMV8pEaGxm802em3RcCt6e9P9pnw+rhPxqq5ixI
0mhcdS3V02JG0Z7khFGRrLLnB9Z9NPiT0heUB5qvQyRlVQ6tsXX5ZEhm1MyAjlzmGTRQYB59C0qP
F17IiWOyXw33RwAfvR011CBejYUjgIMO+LxUljPbU//Rc/57m0vNsXqLa0L53tgMduh1IRpnIN34
7mNs7n015B+rR5qfL44r7FKH8T5cbzgTnObzyrnnX+0S9JI31vOiu782Fr6wbiGWH7M+/+xfyczA
OGEdc7Rjm5iVZZ1kwhtZqJTbZW/KTZl23UZiTjMmVDipdRp0scDlqIG3PgfJ7vNvVMmruXiF1P8r
mnWekm+14xGOiXuR79LMFGg7mcA9xyz59IOnzjjV2jQymW0iJ9C6o1xh9ws1VwokhPJdRhQ52Tup
HhSAP/tvFKxpgB6Hv0V9l1BoQLxvdpRA8SB65ct4OeuWVtreWow6L0eKVULB53+k57ARX84Su/kn
z5oV+I0S8flLqBG5BQ/J7ijO3NCVPWpQxFhY7+e9DxepWpcTPiIFsFYOZpjmeh1JmhHr1MsP1lRV
PjsKnV6zVcyS1oNoKcqMcTIEHMUkx3MpAyy3O3pXddpwEPpK6CY+I8BI021jIwyGiBPCO42GTGZB
bRABxR9DaWyEFVXPQQrNm02TF7qPejtTYRudFNqXxzp2AehBHQUBxAA3jPVefB3zJezaWDnAWE6e
cXfmLdYgkk2cmWmACpaYfofx8y9ILwxBcbQeLht/b48NXS+2HVhuAG1grCuChDo1K9z2BLAx5HOo
+pVnd9O68eXL5SToFKQXaK80oxifxsxtYZhY6oz84toaULRWPN3tKf9jejWqD8Tkm3vCg/MRIKGg
1RCFJhUJJvUaYKdPTpA0XI65RXbQ/iJExJDbfIig78iBDkCgqzCI71dfD5Jbyp+fH/Wb5ik8/Gvv
XQBHuDeqVb/Zqkqpx58H4igJG4CHXL3onujvFyBhCOXEGj4/jbaymUOueehzmou0gnsaZunASj/A
gyuskkR/1WeTxgBg8cXtSo91laS7n0GFJ4ELNHSgpqrlas1DEchQCTFKuXBONg7Vpb5jT3cbwtzm
nGAyd1x9s49kaRsJUqDGXgFIUdHYmu3P9avKUU+xeyGVkv7eQQ71MxWNp6YQIF2cDVgGnurwqVqA
ao04fP/9gvUW1U9A3I/0FeJBuXXeszD52t99IQY+q8TTZjfjx2HXxtszaYgMDA+cAtO4VpzWDNBE
i/kX6w8iPRxO0rPudDP/lb8QRUxcOTaL8SPjYAIWpnv0c1JiHTLt0mph7iHpsYN78vajddPq3/o1
/O3xy/RGv4MRv7Rs97ovyhFuvXbQpDYljBgf0SKhCnn8LuBrG1MWwLdzQeeR456rfylZMggzLNk6
VTceQPeThfzzpz9ErKWLwYwScVHvNw36cnSYljhJ9irP9F/Fi5ItCsrin1bd2cbdZDyQyChsdQl7
7vb9lkFeuQ1BH8Ta1ZN/23YzYdMq4J3zkKrIpza8xU1q65VO1tLqkt1sZKyf6514SXy11JYGAbAA
7GE6c2DvMrFHMFPp2zkA7X3hPykKEfFQtduod4oCLEVFx/1NgvLZFf0NZ9QKvaRgpDqiG+Om53gv
0U/rfXxhQ0ZMca4L37SgsD68JEDBZN5SSDLVPBirkrmKma+3GnStF2BE6NAWBbIlXsKr6rAKvcda
+SyzQz5wdu8IbAQtk5GC2BzbDvaMcLsONG8FB/Hb64E7/mHUTnhf1PKNIpwZOG5pgdTaXfvexYhO
YdiMpLRs5hXTzH9eZ6momGLwGan/jzD8QP4thK7hYr+7/y9fPGCinCSttiLLarAxYJAwWa55WijA
MT9TG1O1MXoYWhICxbe1ozEgPBkI++q+eEOFSNJWmYAL94CoVKYMFg2nvbfdtlQZqGanEbU442Gb
rsnGLEsndSKjLfCZkMW2PQ2xN5uyLY7N5BpqFKuoPMqAD5WbajkTWVd7cgB3XAEhPNLCL7sCKJ2x
OUUp0+p8pNxCb+pyp/04cKbcSDW84EYo0M07ypeCgsrUgZiBSAV/tetjyvg7reTR1W8a3ZZuBnqR
d73PKotzb6xRlF3PPSQ+svAJeIyIprsExAJXpXCqBWIXZIk53Tn9rng96n63/MVBeYRULdNR8fBO
nx/aOy4ZL22OT/MtKcT0nHaG4sdK7e/gMRCKJ9dDvpVvU3mQ7BwLcXJ44vKQ2ZxOsUf+w2YwUPe/
xDV+Kc9DeoB3dsLZjx6+WHnj+E092P35BV3qBg2cNusKUfUlmK0fJqTzC1zW0+ps50t0W1ej6lHb
/+yZ7BDMIbV8UmED6TQ2beP+KppVLED/uOxs20ajKEOpujxBYaGXnRdfevnMQRmKX5Ht8V+Xbr8D
Ln4ErQH/EcBqPGO7NlWR139C7rNrrcD9AKqzWpze52Y0erQUbrxSjImoNkEycPoy8XeA/dbEN8Ah
M9S0xpLSyTwn6MnxwsbTaABXav1ZXjC5zLG4Bro+dIK9vKz5d8WhoCzfbH03US4Hp/NDW/Ymq4B0
+gyqMCg66qfJuzEfJbCE54jUFika9tnGLnhACMP0HZsDCAs81Qf9AmjBLAjHJfLLUYPhkgeVCaGy
1SPCC0ujCwdYKv7aDteHDvC1XIIBQAMJAC1tJtFY2xaT6SxEYupJaDcd6pxYc496kIXjIjx2yczb
AoB1UYivJc4+EXw0iILn2jtdqKdldEv38kFTXA1x7ubNNMRmKGFJRoxfl9Kksb3QB2gO/EjAkM66
Yr+lrl+JSWdIrld9Tl/l6AGAw852dKMFvGqnisRiXV664RqHYZFoXp91K1788cxMeNaIaIpDtU+w
CxH6m162b1HfDsXoWTYKVaIxW+cUhZvye4i9EhNo8xevB07ok0fNMDu1zV2OEd/2hLzr7XNWnLlf
7Cu4un3n6aLph5uFYAbhyu/O3vYYZJR9S2q1lZK3WxZSqkEAHe/lGv/Q0OPcpyLz9aYQ/dk3k+wa
5Z51qjp+qe4eGPR8F9kiqAU6YfJdC0IceztXxFbFVSOcsb5jDM9G8CdF+7P/NABikU1wWRDcjYta
uktCVUxQc49MiAIAgsw+XiuaPZXhNT+jkyanKykZ8U1hoeQkVvFz+27yd6fxLSkCKvEZ9rxBOmSJ
ymPGTerTODC0+EDm/921h8ZXl8R0ir4P7AhHM3WBjeWBNW9mLGCwrDvYLjonneDTiL++RinrESNE
17Ki56AU96rxlIn3f06Mk5cSN685OaXxx/kU/BNeHlj2BW/6dZL6UrOKiVWIaEqVY2nnIu5FOmfX
xXXuBEmSopg/lvxxaNRnUX1FcGIBNkRiMljgt/QXEwzdTr4icZJhPTjQeDyiDV5BjUxRwh8E3uWG
Ig4Mxw0MOnuDWZx2eVlPb0Fnr9vsJbNNVBjVkZHclyEMjjlKK/Cz8PBAmEgGy2GBREXxQirdAuoA
n4p4r4adffcf6wr/fplF7zV/iK9x101DCFCXQqeNlSEWVV5KL/fPX93SNLyVdEnBxOqV/2rYoZrg
BsZTkylZTa2mhmbaoes34ZuGzRaVTeSNcDtj9WELonbsxggSdG/QSqDxlAIN4pJ/Xvk3HazHzmyT
OxfIiYoH0+obYAcTrE5LMn1ixIbeDuS2O13kirx6acUIjZaXx7/wEUxMPPjoBy0y6d7zPaHWIV+R
c96VYiveiom0cLrJ2jdFEWyROI7NwwjQ1HgVQ3FNbpDh9pg1ZhMIrjo3lB5L4Wx+EEh8AKK44nIn
/+RpxWDRoTx+yzZx5RJsl5yeh1XKh+kKBB6n5iUJO5UN1MdgwDLwcaMWOWJJuIeumMCih7XCXMJP
LzXFsiAMWvDgH19A20QN3SWo6zEjxqxso/Wv3Tp+C1Tef+yq/70qYEOwtQuuLRPwMe4iWGf483aW
Tw9dzOPKdqhPzNCDeBWqfbZWgRmw2RUoJJPGddHujZwggAJoZk8w6tlfa5bwyjDutsrYtBDv8hOY
qa/ZSBH0Jlbq/XhGejARCO/qvauEdfF6GLXIKA/iZUpDE+xDRDzQ38SlWv5/y5snFn/uKTaOWp5u
5/Ip8vWLIX6hn0i/jmgSpUh4Z2sf/SeipC3qPH6PpdPHyoO7elcnupzKZ82UUxFXZmEz/ku+aode
Or7jvrButdUUepGAvxlTI0UEbtQ5nscEDAdtPYCrkz6QHiWeTdYBhD2UNl9iy9zYJt/pqx02mLmG
RnxjGgEY5Lgw4cYwn/a4jxvUmfJDXf6NDJM7N1/wFNf4Ak5R57yfrVwpfakZdIzMuMiS5oliLWnU
qsSxQNzQRoo/PUbc8VHVmc7MrPm6JtI2iKdiTAcVMlGLAjalt9HXObiHQC4xCydIFxBLjXukA05w
tnsmVTgTb+p/d0TtK2ZFtJvcwsmjlBHbEik57eu1e7JOTL/XTdPPDYvAxmA95B3PQkIdbIm4z7U0
D4y3X0A7bzNUpTv/q6OfmKx5f8S8Unw54yhQjn/PgTT9JHXNEr5ZFhPNEmAoZUCrVSHvmM6XWLLZ
j6+W7eAylzeAMAqTuKuufq61njQPBtDo4hehszQ8unTGpjfSHbyOVnE3kLPoWDxT/bxuuIFugixU
/lHY/wz2i3WVwFg/A5dcA9GKc3a9bYAEpQweolHHUx4kVAefp+NhSboxLG7sGrm5xQX4DQfvW4Hr
0fFaVarsHVH7Nyhh1N/lyhr4CA+vdqse6pJC5aVHEKld9rHQ6NAmPAa35fvdiDVZAKKaOFDS0u5e
Yuudpj52qiFH1rcj7eNF5a8NiBOXsogNx3KKOT0spLdJ8oynZLzWFtacclIL/vrblY8jzJlKPQkc
zsvPXEve7QntuU75Q0bRWrZg/SdrtO2FPaLyhaCIPoWwYruuieJlBQ76wV3eaUaqUSxzN+BW4jXS
d78ck4rmi3C4uRAHnU6xrMxlod+5UmnMs5ffsNfBpY7n+10s6oAIYcNizSMqUzfSi/J1mge0sc66
t/w5KV7B2J4eLQQkUecYkBXSn1c8JbM12lU/lyNg/yV4+8BBhiTU6bACLvX8k50tMHjUgp0WfnXo
ZG/6E6i30URoYU6gAH0n42qo7kvYqpGUDMSYfiHy9nGFflg8MPv3k/q8h4VKxFJTiqzcGNgLEAPE
GOS5jSNycb3EolP2eahnb692D67s9dh7/fZ4DtV3chYMrSakyDwNcLnZyTFHlZkFDtUgwenySK6Y
Odvap9A80mI7yNqCvRSRK6qsW9XO3quJoPKHdQiZa7uK1mTXdF/3cH4WLvrDBBKvj2lI1f1TMSlA
x1JDA/LWLJ45KHnedkndqc5zrDMzlN+zFf539U8sf6FSkMnCQxBrHpMbak2Jw6KQ2RgP0uSEbXp3
AKeILG2t6BVpoTHp3xeNm79boINxQ2AetwA91l4DZ6Ugx0pv+FCpUzJv+QoMcTKsj2GSRtFUg3KX
81scvU2TtNRi542xD3wtDq3MILV60MhxW7EWZz/heu4TzuvNogItfEpAWol3NUmPHHyBX7OxzJbb
WaqGlbJBQdti6JwYta24vgCdM8VJCVRt2FAr9viXhcL8OL6LGyDqR6xP5cHzFs9nB3yOHoKjZdFH
tOO+046mXKlEiN05+tVkVubCTOepPRcfls1kOPQNMQGN85hu1YVFlUqSpy/C7rJ1xWOW8W20vaQd
awNQdrTXOEJfVdj7cberTTYHvshPsQkH5knpz45nZ2I+Xy/Wa9V+YXN3rSTWqdx9THT8oma4Y4ED
xAaOViL0kCShs8yxGd1E5FfrpjBUFRP3SfED0edh5wkqUk/tUaaxu68lNVgedrOlG4MvCOVzpOQW
Ln+gpGr5JtcdFtcEdsdorLiW3xvv4rslsazxVfqF5lla8KV8J7okSDIGk5ASzOZErHLNQmHL8gTb
zP0H3JJal/SGt+MUC4v+1Lq0uWg6ip1zw8LKjuEi8bBIrlBVD8uS9rm9hl3BqJ6Mr8+b57aB2tzP
yNjQG8kOzUBaT0D0QXe+/CujPj3FGP46LqNwMMUvrnan5wxzeBM2TxZJq96Z8aJT1EqfNPNFnrDl
JcIT0OqTmDgJ3shSKHyuqjW9sfiCDwCs21JAXgzUs2KEAct1I9PfAjU/be1lPg+nfAqCt0RCaBHR
SHnuozXk2cZN9LP+SnSVrolexc3V1QRW5qtOBzCj/ByqY/eJLloC4yIYIGN6I5BpLVmzNm/s26rO
RrAjzQ+iYha+Kcyw5haY3owrp6IKzvoMRtFNmrYruLm0+6dwX8fOS7b9ZaSfsM3XJOrKkOMwza6J
N9m8d0/5dXWNPt4PFX5jWjABjy5to6T9azOBQhn2+AWpEtJKlPf5UnQUXygW+f/AuWHGPuaUbYmE
T89NGp6+xRogJJcmr2umk6NXmJ5JDKHBiwmablbg5OntAA8DGMWTBXAJHfSpED11hBnkBPsZMDQ2
WRCIK8cvwoM+1QfS4AXZA6mU1ehLQf85MNhYpHupcV+GJXjqec+UPoD1gr5FiCQ9LhQRydKYiY0b
gA9Bc+5Nzx2hx1407lsvAaKcNw+IlTwlXcrKn29o0wQy9MhVyXx1Ijqg9QIf3WRO2UI6cWw5XaMR
HK4v+BVQbFRPXCb/LI6KtNr6YpbUFMAo1x8GfMVwK4wpweVhBa4g+SJu1vsVvAVW+MnrsZoDB+6C
CgCrx3Ms0ApTV5HcR8j9oUjof8/PkjbqkW5k1TCtCRmfAA3/9iZ+rs7us8lnkiI79AeGtp+bPMf4
HaBi8tKGCwybMuId1taOUKcTN7p+X972f7VyVjEp6TPpICnBc/PR1e1oQP+nMWNCyXY2tmjc1NxD
yZYO1/v3K2u5FursS7lEp90H4rNS00TPgFVehiE/1u0Vwxe+7IES60SYGIDOPXeZvfVJBI4US+Af
jeXbOzG9V02zV9f+cy5tFOJiLhGAAdlAk/bt9xJgVTPnGL8cX/IDCnOvEex9HorH/TgDcaa9dzM8
KZjf3JNf7ZfzXy4rV5z3raB7oIaKkMJblScc+l/dbfSCNXPIrArHFbOiPiVcMUq2a28xbLIMo3ye
wHNc8DxhORNcbqMQJ3aIFdDgqOwjHxZD7ApiMAHRco7/0YMqt8eU8IdHDu7AcIFkXIXLAPBxofsy
hqYuy3y2//APPJerqiAKUqCPBxm3TsArTUbFuM8/wl2iWYyZbtRImb6FiRZRJdpNmNINFD03qrFE
J3F2jsUt7MIPFIJsEo5kYMDjzT4KmsiHXsqCtW8tRB7vdxTq6ryCILAv6E0PDg9mcwSq9pRi7oc6
1cfNSTtYbJM4m0ZP1QSESofqDs2bYGr1u4Z0ZS5s6P43q1nqtAvDMsEq6i7HNm8AHd/Qcl+hC9E/
UBRRJkG3kIYY4Q6UZK+6UW69V2Yg1ezpgB2OUJEK6dYTZA46yEHpEvvhNK7bTyhrNWx8afVresdC
u3q6Yb9c/G6RNOh5TnhJoCLWBr4MJl6vk+tZX4ydhGln0AY1F26um7dn8qcBIrVXgS0VnnG0JIdy
haicwa3O4lfSG4M6IV3PfclbSSZqDVGLVfnPUji+2ePtKTMnPF3jYpXJvGmPHPiWP0DhhLpj+OLj
mEVYiTfzTSr85DJ8h56Po9eVvdzOpoKYZ00irQzYGMJaTnz06R3RrxaXmK/8JHUJxxI8k5dq74Bl
WKsWaGhbZjJvraMDSZbBMXzTlpV4R0WNYR3F2VJfrQ8jBXh/RGTfbS/jam7/hOdnbcug5dPtaO6B
dqLLPCZRBByWfFeODUWljpUEULRZMguwpnJ+oxiSA67bF9yVPVxyUo5AOczv5w75fwp3bIww/ErC
LP6rMpBPHm44KlOIL3rNmJajC0C6su31bsYXWLiQR21NmYFmskbpX8mNVw31Uqf0YqKKlYhPLwwE
r7CLUsDygljzuxDT+0yr/me7I2aPg16eFKdkK1lAmdl53nIygKPTY0JUoN8IexzUYcOrGxgsIr2S
d9XX0AUnGR9nP0ZnmSNzAiNn64jDh+9p8U2W9PAXlSnGIbxWxSw7QfaklDvEi21ZZQFqqnWVjW88
EDYlHJ291zhIJMImjZu+svT7DIR+y+SN0FUd06hSfejIE2EyKfJLI8lqPKk82JfK3YHUeGBs9eBC
vlZpsM3bIXpFIhY5AzaFI5O8BVD4YmQ3rCV4AA2Wdp076gFtH5B8KSD/KFvJLV7WljpgY/dbLiPi
uK8idJxKK4ULjZv2ntW6Cx+Ezj3g0wXPO2clwpg1ehRK6rBFQ9P4ADILDKp427tfukkOjHHbNqKb
2tLWLhyZIIUNWYsB+cUphm0vGxh4pjSbC/ccGSi41XjwuL7B3cXvDROhBxP5ezSpvpZHfdqwrok6
GfKrOh5BEIYQz7DqWzi5G0YwUJiN8fotGdpWWqDa+sv2XohcgDN1ZrRcPSpEHxKoaYfALFNW1MRT
POeDt1IfQ7X1Wbktacy3bJBTov8GvbLXlfXprlnszUSuw4zlqdedzHuqmCKz8STEj8cgW9mICwIQ
fm14Vhcz2ZegzOKpNTtwugGN7meo5oJY0yqsmTeJypHHDNaLzbNb+ZA0ky5wTe3rw82gg+F7Gskz
OGAGIoveOgVwrrjZOLXVDsVBAYr3U68XzfIudct7/9y5cRG5D2aZ9qxtRlGk0M3KWjreGHR5djGB
3mAytkaRimg/29ljYjZRSaFVNdIt7tFaw05wmicmphapN76J61sTPx3oe2mZwhnHlJjbSM/yu73O
4nd9acAy0EpRFJnzb+7TayTSp+Vzg3wE/mo19NU+RPItM/HpzYISnzZXPCSuqEwH4czZlCFR3VLg
6hmCR8A36Fi9X9VoV2SkSR8wYw1O1jygHE9Pkinxi9BdXSG7+mvTC+9cl5FVwcnVNoUQEfb2Ew+g
kDdT1gzmlOCQhhPKqSOvsaP/6RXHGGz/mVYkEONwXHpgIv+KQ63INardVhlQbAuGhZOeG6BrZFlL
Zgcgw9xdyN/x3xGFiFW7OkOqB3YbD+eEW7J6qiL/UA6LWwb5Pvv5MIDsTc5/VV0FWYhcaMjGJYTH
QH3nhFP/RsNnCnJYa6JCW+xS+ePYARq7JFGBYCUS+0EOUect4Ceeimm6T+LL0SHx2ZmxuB2dvBFc
pt3L6/HGWSfgQPXtRLoiotaTzgfwLjTNgB3IJxrjhMFdul0C1iF5v9mWl/42N6t3DhXEY823T+bY
zuBkRXFLTj9QNt5hb8Xf7gdWmJZ7QMobGx0lbFXMtS3ibuIY7ptFeUe8SMURBZbTyjrhFrC3U4BM
OnZdU4+gCRelfpPLBwTrTWIjvmFEDAWvSJHBzHqVz9fw/t6FhmqWIKnAJ8qSSsmiDOHWn3trZ/r6
ved/GhBvomf5bVIDdN4RDmuPIuC4nlQveLEArITWmE8YNTa0gzp9oDj0Qv0tj9txZvUs4cTS3xVs
A35S+76bdnN9NVzl34LKQm2qImS6fX+JUHt2RX1CcDpF8T4D161qyXvm0K7x2IS02/IuuG1OwNvZ
kUUUqb/ay23XHBxSRi1QPQz8VX7fsKtf0qu6OTPQpyWv2fd6bZoQmpQnkLweH/T4eUq4/bRXI1S9
GRUBh7nTNL7QjRnLIEcOsknDIV5wW9yl2Yr4SelDUk02RdDE8Jkt3Fbd9M85YL8C0MXZ19KY/Os+
aaahsTXtFSAZvyUgZSFO3/HcwVc1vTOylQzGugpktyeMF8bkL0dSNccOj0Y4xvm7DCKyNMpu5+Ti
qZdH2q3DX2mt3awf1l12DpXOMLi1BOJZQylfcdyA1cW8nKlpX26e3IAL9uAdJHG9QvNpDF5alKes
Xag5wsEHU2OgwFQfiqi3LdXx++52uOB2wY7Lub83u00OFGFsUDHNOE/ROBtmV2cl2VB+YxaSgKGM
ieWQBDVsplwHLjshC0l3+az63xUYaIqKABED3dPK1XBKft8LXqJ1+leGBVfNZUJYdzOwUregJ7jP
IRSweR9qD6W4ZcF/T+eo6gMUDUBFNVocIJzL5amWgWr5fQtb2eIi93cDtnhgPDumISSTw2mYqU0R
tmdo+1GFhtfvJK7KCY+Sazjd97VsGTdw28lS0bkIjt+Jarjr6ru4gOVdGt3ltAoSB/17c8ux6Eaa
ETpdGT0/u3WqVWVFint/TwOyjv462YVuCoRupbaX572GF25C/5OEy3n15wggMhjH1NiSORIDUH2F
J/pCKqAb4gNmOlgPTMipXFCKlMcdGFhnWZ38LuhmSEQ0QzV1ACP1OuM6cat3kRN0D3ApO5wGlE7b
sfit9DCFxGg6rci2ksZ6inczpAnHBv/atrGk2fAnHzS6sH5V+zDL2G0WC/of2j/NK2YYydp/HsrN
zUJtTdo6Ec+JpLvfnSP+gakTh1knR57Bwlbwl9K7AAvDGSlJtSrFraQCZerbhEfyc04c5gYkjYaW
uJYjvNQrW9fSM41qpt+Ij5a+jJ0ttHINgTAWOV4ZrJFRwO1ISz2SDnbT/IR24Iau7y/guXGO2NN8
fyimMBQoiGeazA5VMO6PpDULB6OwIr/bvnGkuxQRe7lOgF1Hekmi0xc/4Me8km9EOPNJQAP6m5IG
V8ue/zMBdiJU29HYV5eJS63pdD7Xq4uW0TQJCYECsrrFHGrZDKsUrLnRiJV4xaeGrz6s1O+wYhUV
80K5z6BJd31QgRMxKCur6IQNJqsjxxs813YOQ4t3B0UrjwPrk7ZARVIzTKbDXqN9ioBwXJ8hfwTx
x1yLkkJqA/FEsrhyAACg++KQA/Vp+MqfTCxL/iagD0R4LQEXuQu5K9LEwskdTgu4zOCXlzWzqF/5
s6qx239DGfVfh0YuLjGkdgYIwzimG1DtnBcf1cJJfQDsPV61dgToFdXDddTU1ndTwaea9ETrLp0A
oBYqrf42SqPG773rEHI+P3fgGaLM8PAPLFgosnyL/lvHePZXzNytqr3+TQD6moAXB0C4zu0PpFms
uVoR+Pwe7HAe+gPyBkJhYx50lKCTUN8hkQPeYCD0oUlpQ6XPTpZEi58mzeRucRFzV5Oa6XW0M1TC
/qpNHOyWig02+4B5Gq2lxp04cwJOQqcZqAlV2CgPZMLF2KYwwcDxPHm6VaJskhxas/HjlV3WFQsz
BKQZgx7qo464/UwsYhc3RSAf1NENRYrQs6quXLGqD7qScrocTDiZXFPqy093sFafOrr+L+htBi/8
BWrsX4bg8ABBYQlYh/Dbb4FW0ZvU9crIYHHkT4IOq1IqGn2nFn+8Vl+sOXSbALCvua2byAalvTQL
h6S+xFm9ObWdhssFtukJxvkdJ8CAGYnLC8AAw3VRkD+u2ko/qbEdoZhOCZfNcsmto4XQluqoBeeg
Q/xJnEptZnZHw+JGBWxSr8EdBcnFW59cP7Cm41tgyxmdZqR45N6NcRGfUA3zqHS/hmX7f/TRYifs
vyAhCEouSi1a/ZP+OfYMuxmzQjCDuC4R0vMZkwCLEQB9ONhBsOXb5aUOVKuUWg6iaL7llU/JnvSs
kzyh2m3m4n049u69/4NlAPK5mzf51jPv2Yurnz9Iz2O5UBRNk0+j50JGlyqilUPSfdixu4z9SGy2
xUDhSUPGvTodgMEadpSjnHKh4+TSP7dqxNmA8Xry5IBExtgxC8UsdOajmgb9doOZrZkd1NDpJkga
y9fbRPRUMSfE86AZ+6U+MUZRvl9iTbSu1lVyh/fm9Run75GXgHhNUAYQF89XpV4yxDl9+eUtbffY
WVHb335yIVPQX2tlUjok/Dtj85KlMlfCP2znUyt5+llfOCU4M/TLeRSFPajbBGHSuJ+Az6z9usGy
73z4N1a80SCn5gweRhPOfnJIgZXPeYYkTmQDSUeoQoHbUHRZspmfJYKJhmvE4t9T9I1ARODWFyd9
8qQE8GRsDtVaJaAB3z4VRC8q4Ov8/icQJlMHNbtgo2t/edhvQqS+6UBjNSwDe5CMwnyodILCHneQ
Lj12WgcZOCva07qAwNYSz3GjFY0fpd6zMaHFWO33uIQYQ/fyVP5Ejd0PP4F1SMev8lnXOECvhF9v
y06H3wnj8aNWMOqD71F0hKL1KVLRKCLvBlZjpIbjd7bNc76PPSHpOINPrC6m5qx1sNV97o6I0hxS
FxRet/0XP4k7kNFZhCeHZ7j4v+pJLNDn41C31f1k8e6ms45XoQcdYAuZBH37h726E8iZjBGDQdmP
yyC0NNg8kN2s7oeNyCIoacL2x8WVdJe1j9TK0r5R+oTYbaRShhkiD+6OSDpsZnd0xhbo18x8q5O2
/2G+7PfKgIBLNRV3ChUvBb0erBEwXVbFTNgMQYt5dqN0F3X2VCtLZYerUKhjJa8dgvcKvzbcQhBB
cUsd3CcuM+nU6N4AtAYmftfyZpDLAzTedurOmGFxmj5dkuDLb8bJMH2Ys3xX7UZjE0K0FWDC191v
ocEOY5vUMSKC2HuKwMOJidHixL7Ip+01dt95pstTwK011vPDcxpfxetBys20Jl+nSeSIL/kZYgIS
TN86vK/pIW9RQ0yvHQUwRkpq7vuT/QYJK8V3OaTyc9Tn+9rwDxN/vGkXTZCoT7tOEMq1t38HB4An
XqhVruL3WdFowlheCBGeA2JggO4h0FHWia8IiYGqW8JxOUIaOrT9jU4+9DvqI7gHyeTNwvP8dcqS
EuEO6BRVVI36ottZapCmGZ9t4MflWKQfaMAFA2GA8EFnZEgSPqaqe+PG74nkESZmb+seqOJArsi3
Fbp9RxagW14IvS6y9guT61HHl5eaOKqdo/tOVy8nYL35kob5lRd15gR+oxW16NYDn5yewuDEvcWy
9oPP+H7L5pH2KpLBAoN+DGpFWPre2Hyb+Kmq+CSeCEYYbTyPGOyAlgaARUU3wbU677DK0nTACI0n
xh0FZ+gMTHfAG/2NU7mtNDATYk1wUGSJVadH6R+Ptfd06Q0g3H1Sj6WN59pN1/EVPGj5r7nsXqVm
d3RkhqKNBtcoShBWoY0YEGg+uCiIYJyxlfp0tFVlddZpL8yY8mLZx9WISB1e1Bt02Znwc5fbBzh/
dC4LT7h45HQRXBRnIJL8yrY/MGtMFQdOvmcMmMQQgV4JQFLYGAKD77ZaOlL0p9bcj4wcCmVqXWUa
8ZsRZXtG56rsUTJk3yl5wuZVHW1zV7U98QtmBiIdIDvyKCo9G18DhnVtai7qqYS/KqFjC6fUhMMW
wUsVlx2OaFZKypmcuLYkHDknZ9Ii7uXvkBtNEcW+39FIR7/SttSnibnymhRbAd2K/vEOoZfA831q
BOjja2de/uDNB5IaB/I2jVikZRfhq0q+itq7e314LtzFuttgoYmHGlaA1A+HJIQM8KtCYuSmvtjO
n3y/1+1juqghwGOZIk6fSdCuzVXhmxq2DnZS5oz58hwDBGT8Er+zC6jwp4ILI8Pi3bIxyB3lWDGx
/3KGYlTfSP4CW2Fo1KxCy808OCrwa+erMWOHiCD6tVxSw8R8nIopxtkwjy0rS9izklSL1I6u+T1i
30Fb9Lnxalf+o90+nn3O+ffDeV51UjijJbzHFn+hZQFS6f8h75CrdtI3Zp5OXabMcFJawpWpNK6F
gbVkozkIVe8+760PGEjhAxE0S4VutMQP3XvMSobHiWNY065Nn+tI8LYecYaHSIL280hknW9GZCwB
0C+cbTqkXucM6HWU2PCQalW6/2UbD4ZQShv+VGLOB4JzGciBLXc2KPmdtK0vlWc9z32h+NNekTbj
9SHBpuekJ555lZZKfLeY43gvM6qgXw996v5mf2CoLAGF9D22XiET0+5iFmorYUHozcxxTCsb9sUo
h5I12jWko1w5AKEXQs00DK/Gkgbdqob+FoieklUPP2p6+EY49SLXvBgHVlRUTt3fBGr8VBtKnzm+
uf9yqutN/vwuf8Clj/oracrr1IkPyVgyU/ljP546h1bN/tP03L9h3rinJUK+GXG7gFkpXYUu7Tg6
CC0Zt3PgvateKRqRigxPkDVMASR4N19rJNxC5I+zwETA51swN/KpzAxtNYkNetg2vdHcE60CLe1u
YJzthQDrFnJqeBpoSykznOm+1l81fRCbbBDooRY1AB+L09FA3zjbNbPw3jPfBSroWRFTy5tNTIZp
qkCieB7M/6U2jHUcicbcyfBXzX7961cFbyIT6zJSobQOWWlbLWSPuGJOzVx7EzWCJ/h1HDQwCdDG
aD14AiwA7yVraul0iovWphYY/r4nWJEiVLMfvG/YiIJEQiuaSO0XBXdkuEd88Nu8JgbHxcVgV4No
FL7GIbR/fDdFAf76xf1N2xwLamLCuy5C7qn7fKWANAb32bBxeaw2oSx4YkG9Jy4vgL6iz0z78f59
vA8eXcuF6c9WID0V6EvS0f68U7ZIIWyiHq5y7Vjmg3C2F8oBfZ67+r59QvHpA3LVQE/waKZzWIVO
epzfcwBopXW6ubh9yq1OKs1ulCiv57akFCLBGj9d45oSnt5QAiBDiTEyekhP0FX9hftjb9d9K4mp
7gDjNbr4IK8D9WJhnhKFqKN5nZqVzvAp5u0MC6HhUhQudcDKGU08ESZBTWzYZIpUXr+vhfxcSQ2O
bm+Mhu+nhHJH+PyTGnqKX1jsNhtWbRLdUMi8/Lka7d5gCHV19TfKDPycbQJGR5I8NC78hJD5yod1
vmL7/oDP4nGt0yTV7mdY8SzK5WebBsSOnJtQTy8fT/d5Nu+wg+9SRwr21Ao2CyUE63eewHzyHT7A
GHsggKGG1NKHA0ct0evhXmJXmE5i8dkxNykZ4YDe1JfdxXdGdK79k2HKO0GrKhtAME9X/OkiDCbu
lyo8BhgTmAeAI0yv9BdVb7bBuYwzQiqVNBeo2epVT2SqDLhdBhjZWI0AmruPOhvZ1lKPPoSx0g4N
2XHtk9gLzBwnQPxW+7TXrQlwyJ9VCjODUgkzm2NXa7cVBelkmHqPvAc9dhfj9vFR2hCCRZqHZLT2
QZnquvNWI6HKfPU0lDJGmfZcJUZea9X30zv4AWzZrarSSAIf49jZCsmcFIj6bNKIut8ZFeX6LOvl
DIsoZJxZ88FZH1/UFcGU1vL4wNCpX3ZOyyuW/hdieqkOFAL+03f4nrLwu7c7nGdkMIA/brV6wadY
srwtL8/smKw2gH/7XY/tlZ6MFskeOWbTkJCkVIfkyWk1mwZqttztPc0NQ08Kmi8ZhsSQbrExVW+r
jXj10wYcuBjHi548mvdDM5m2SL+iz3uQhjlgAEhlXUG2Ubl3SV8cJ7NL/C8OERHoty0DczSxEMdI
TpRNI5ipT+hRJX6GHa+LvtnNAnPDbODfRhS4IXC2IUhJvKjM1CZpIk/ijq+VzrqO0H5roQSSPznS
NchBR78BLCtLlauc1sfMKJZFAhS5kw7a2zzU0QXm2Kxzg++wEe40pFnsUMI/zSZSSm3S/K9wkucJ
i4v4asqo0J/V+WRb7yzlQ57w8ArVIhd9SUFm8IsxXxoRQ7yiDZEdBy2eqsZE/iVVl7/DPj2ggK/i
0/QYrPnJ9I6H03I3cs0JNr7yICkE5xffzb77Q+mIW01mu6JGEHI5BoBX2l7qzqcV/pTCspbm2HeR
Fkv9+xjyA3eRjuZ1KyjeLuWJopiCM2HmfrH9tfiQ11Zr8gpudpSOkUzz28uqo9OnSP7Uhv8zQ/4w
rYHKe45QIecuWQmFjd75HyQ2u0bK3Js2wCmJlhvzXVQJOouWAVzt0TNWUDZgy8czZkp06hQpTAyL
YEIEIdWLdO/NOHnM9WWu1j74JZ17s6S2hjkK2eWPC5WzKzVlP2cjEcJ+jaDwSXhgj7pjkG0HIKDH
Ro4BCF6Hx/tHhNsEbVQshHMRAKtuCG9wt3gPLFYqPfFFw9RK5u2ToIdGmu1TlfznE9/hyaAp17+p
OcyMxQiC7bIV66+81RFuSI1/ymgd5uaZ0N1FFT3KFPIAhUEzJ/xgsE2ZbGXKK6YrqDZFiRPGJHov
hROJN55nJmjoSFMAQcPxq2tKIQor6UdVGP5JayCd0kj2ozMGRyxuGnCPTsvp9L+r9Nm9LyjUcBlr
BZ1kop6xnIPwE0ngtU+qnA/7Wj7VhPSVYRAptoVPzHaQJw312ygMRB6ag4ekn2zgaZ7XflnpQWZP
NZ7lcLquWwMUqBgmLw4rFnKIjRTN5SkUjtoJpkV6Du43f+PDRdJbPv50xL38bcIFinPWYKECFg7Z
s5aPcq5/R82p7LfQbM256QQ38ndqEaMfbN1UPd4QTfNyjGPwR705ltRAzRITxTB+IXnbvPUW2E46
kTdGccOBAdL2BiS0KXO9bXVIDds6oXDhP5DA/tn2bYpTRJbm2pw7cOOmg9LUU/khwXNcG+obqjxd
WJEOvPxJr6TzQehsyqcZ0PeSgTNIunNJYQTA+XkgU8j1vXkoSR3I5bF7rf+N+G2qRtk2nEgw673h
udVpatf6ulL72UZkJ1j90jcxJUSWyl42jmgm7bfUh14ZgxTNC86CNFuKyxQTb47qh0aPj4N2PgMa
IvgH63LlFBauk4JF2fQldMxoVAC3u922p+S0Y6JrWNQ6pcv0EfkzCjEUUeaKYYaTHNhZP/UshKUl
pdmtt3OLPm6foMArhcWVNTf+zyWLePaPMhBwq1s/hzJkQh+pQzZb2OqVl7GnUSHHTAoIgvmHuEJw
0XeZMcFJbql75aIe0HCmxq4jhulNtHP0keXqXEd/7n9Mj2Fvq7zQFZSoQcJzoQEbjD2ko/7kMHgi
yKeHyi9HB06cHj8zVxAYVIkYV0CKgka7PxX5oSGNflnhr+omzypK2r6Gu+dZnJ8TdIb+lEJm+zFr
Hm4QQpQisLwJ17B559YTqPFQneO99IYaU+KecK8LgZBjcstz+r7ynTPirA9cxWn8gNb+FmMobZhN
BczTlY982PiCeVyqntEupDi02aYJLHJ4XyYexobkz6A4NKnR2c5DKorXdo4Ww1nqNy8Z4yFrS+pL
UHsl12LFDg7+PGJ8N9wPSbyaUjd7SVl0tDzkxZl1rj8uwcjAQYK9xysqcGkYzkHqBeXcbTFpOOc1
nEOCYmFO8q6djh8g1fJ1hAaNGYYkYRmAZYNn7ra03sNTEXf9Jok/o1kdnnouHvtGKp2GkKfmPlkO
BL8xjuzYMlwjlgnucgtXZ6Rdjan0omsYhFnuXNsHLt2d+rAUE1NkWN8C3aFQ3+JBOzM1Gu/dHk5M
6D+AO4EHa2cruOVOyNYmXW1bxjFah/qlpvFtkTrK0tD3q8u5xpyFDEGMaw9yIlSFXvRoOr0Rvscy
JKG/iJ2Vi6CfK1Z2bDQKhfyFzOoUa4CZFii4PedBLJEMtc4B5MzIGWXcOZBfXPkkQKrZ3lYQkXNY
W/RJgV4w/3woyZ+4gieZOWozODwtS7CurDoES1cd3Eouj1FBpyrVMT3wHlWqxE66jn/tQD6g0cAO
ofrhWB1Jo6X5zmBBdV+7TfNMu/T2OD8Q7JcEnCWXHBfhPkrROrJZBocOc75ff8Zm1OMkwQdo/nJE
Ny4pz4s4vHKj6x5ynyqPR//kHSyHfnYbNVuDDat57eipLn2o2MWW735PbtXQrg+ONVfkqwhZ/QJM
mBeNzNRqEuai+JVIavbRPswMbHkg7sgTKrrlKB0APRB1BhPkVAKqSr1HAwEAoU8NpjzRoPiwjCpG
nWExrxKuE+Igec6In5GDGLMOfm8xYFomZTog6fGcVX5FHuTSayQfVrxuRRj+1qUerbzcKlZGlWWX
wZOOVAiY7AejGoQVhRK31mbj7aok7xED2z3+1JfGH6Htsd41gZYkrt+jnu06TCcH73feCDLJPun+
VqzXg9Pd7LioqwvmOTeLt9UA8N2OAUxdAgpknNq0Bkx/hGqFzfOoLp9ZdnsynJUSoxe9Bw1qzue8
gg8lLwESDsSSjH/Ehj8ZFUvNp2pWHcG3kMg+h+TkP4LUkcFQBxZ5GAaPfKf4yB5lSAknId4ZjXF2
lrYZvc8SkaPNF7HK/DfN3VJTr82L19YtO5czq5NKgHYZjEj1RB10gYohE3vTwddPsvKBItryVel3
5T/1tKRWcKcvZvbhCe+wxyViuTW9OLNCjd6H+9/EwzCwnUToga9CdAD1gHM3oBCsiw0RoUSz76uK
ZF6OZjaxWhWTArLtmRNFTW9Z1S4oYdgZaUcavNlldM01a8Lr1VMSbEveXacW2usfE4hhzJ38apsA
sOpFUhyL4Jvva5khA5astL2SyC7DJnIMeuKIy+rK2Xgh/QGC47JQqLcyLWDTa+Ogp1R2UlOHb+DL
eTsHAEuLEwak7Tjdf8rZFddVcloUNsgCgucrO1D2oczkUZNWIhBrTNLR9EHs5a9XGdWMrfJaqDKE
6KC/UNDu3fkD7/WjeswpOxXg0yBO6eTiOcudPgFCf14nJmASsCNeEb2prTlzwU2GliQGHV5r26vC
WywizGnIlfk1s3mL5lUCz0rv/RPFUs2cnBJVMMUalSHYgaZNje7OWlIcz41ZWjTr0LCbBK3EQX25
/ERqBbf1cXEdPvoUeb9eF/sytZaCr8OH82PZYVTW+aD7rTmR0P9sjPm+6OrZMp8umO6Ngn5runt9
dbev7NKDzNHJEnJEAS/PgWbfO1MH88s5I6q+e8GNbS3SPVgPnLErbWzTihmU04eGnxejxLJyltMB
fPGSFw9zdAAceudTQTDmseKLU7GRU6cY/7g7iGF+Au13wxwnHXexSwugGUjXeYvkLyv3+OaX6Ux8
Tb8bWzLdZ4birfjDTEuxSzQPHcaKqmZmyuV9mDx+HTsnY4mAFoe9/fPY0gC7YkRDcZnXddJ1nCKF
UiQZHWbaXtTcMm/8jFpvgv/joa4sN5I6DbMsU+MYg9MX/pZsqbJ/LHfdE6LpN2VHBCkes4F2uhJ3
u5ECCk1sUa5KryZx9iAsmKIWK5y15MtPbWjOZMF5S/WCX6Qr1qsWmloJbk0KksRysmw7+49k2gQ5
InR1aQ5RT/Z+z6qMqaUIbimXRGqSw7La40h6taEbS5LeRHvBkKhRi+lzvIkLg2yr36cGExMzuCw7
Z/ZZlI/LNLxhTgHtdriaFGWkj5E3TS0TENMkNA8iIwQxcJtvcubmlcbGl9tW9RVQquk4KKpx1Tca
8qobChe0MZfK50w4t6F5qNffkoQq7xhD16v1Vu/MmB/tDWx32SX8/dZLpXSgy91GtBL3KhS5tcuW
IiuOcJAPD6l5GLkRkfPkfiDSbC5ICJpqmpWb6EQEu74o1p+gFIIcGjKws98C6LbG+0uNsLDIG/6l
ThcZHKBCBzOpGuvg1JImtCLcx8plXLXhlnujtv6J/02GOi0iCuiVDgUFuOymN0CHe4G4cpGsMXeZ
8g9MbdpdOJn/6NRhaGcU8CX0YFHCOwZtoLIocFdwDDFX45hff0x4jvrwL/qoCWSEDnFDzYOyY4G6
1dXRM8B9THB4gCpP1acHpQcwc7tIUN3i3nK4NkrpkdbIMbiI+JWZf6e+qkGzt8V9+6kp1orJcgBe
hlj/zia27ec1HHcHY3laSJIB7WsixfKLxzVCkunn8wtuFSCKt8BTRqNOWIR98dzstm8WoJ58Vhbn
kZjQuy2HHgi5XQgqHVw9K9bBziBmiKZ0VKpSevQhzkaQ3wee6gf8Dd+Tkslr4UeyMFE5dFFUkvp6
H2Owxl9tL0IrjZlCIJ28dj/cxB+g2dl67TQKz1rX6X3SMIFplURfv94AJBnnhohh4r38o+rFOLK1
bDXO6XCyOPLahRPspyQG/M2YdWp6oNzCHHewNWOzhidWMqUUpSWDtOIKE6VlhbxxzMMkr2lyg0JG
8PwBuPXOxU7zJ6tIXjqdRHUEXd5FRV22m4ncJghClcerjANJ8vLcvAP6HYWN/EsW9ZAMdDGojyEl
TrbbBtlJdzEG6JVKK5ywrMYjhbe/46vWqc2QE1fFinViepEfVrwZ+X22YU1J20kTDlubykgek9zV
0WQJIgwkAFxCOLhfR2cfDbvKMOVH+tzrYYxgIJm9XwPaGt/FDjaPiNKE/3wy6r4f5oMv/XlGJEaE
ecwBlPV1LPkbtNKmv1gyEBdSsoFKvYKgs75CnBFVyn1y/4snofmADkLRrEPYJCBr9ymZdIF2jKa0
X/60o2/Sn/TFh5hw6YG6JKCZVLtpMK8LYIqph3WzWG6fau5j7aNjMM1Q86FVafAiWSCQ7AWTRfis
/rfSKyr/l2eKW41LbCNSeQe7OBqnvcdnPMCE/MBrJOc6sBoEfbNUvZCO39XuULHAum7mLFl0tjjG
pr2EXwG1EU38xgoQuN8BGOZBiQlc5hNtmST/kPNEc3pJogga+M7u2NJJL3cMHaNcSgvHzlPeRCPF
ByyrWhY/auiwGM2VRjxDZMtM+xsro7Y4U+JPNwuyp0Yc4so1rx5W0Ud9JGO246NDr3HXwxof5yUH
eRYpAnnoJXKNms3nyD+r6fUYJCM9DDdDlfRVp2+0MmuAYQksJBLoc6lCLrS6XOsT6yvXunrp5LIU
Nlk2HKPrOtNtLI1wYYojSxxtSzgA34WlRqPxsDO3fxnz3RiyTOWyb5uiGieqRye+TJv0xwZsM+vG
MmGo0sk=
`protect end_protected
